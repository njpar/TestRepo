`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
k1TNL46COhbmajA5SKRiGL/yY/l+mDLK/tFf+4A3HrKrF54pGquF9pt8iogqr6NpcWrTvB/+5+em
uF3qey4pJA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OcMMrdACL1+XI9+3IL77pujXvR340n8QPsMSnO/2DpRK4Y9zF/C2zMEaC+5uxqsE6PwKLSXPzeF/
IC1kWxHQKxI5mk2ZeBSsrFRL5K9uiEjOODHu7ANYk0PEpzAPBj1oKaATyTeE1h2WCQ+08zWbU4+4
//x5NvPGnOmpf3Muz54=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
yV1s5CuLMOTxnsxqCKPOQeVbUNk8NcuwNdhjTikrBhAkcDuYIGXojoKVM+imIaAyGHiEACHH6Ps7
oi+WoWuplClfWkapYIy28TfkKVI83ukfoc02JKrT3c1GPd70i2IloCqFd4haKR3hnMiebSM4p4mV
fkcbl78dOs6wMTFZtFNIjdrHIBtoo1U9d2Cd8VkSvfGTteK2f8lZgZiLr0tbK2PDiYnEw7Pm6dAR
R7whxJbvmKup9gGUlFk8r9WhkRZEpVmmcBCP1wXsYZ9Gbq7tZidIcrjOV0id6d1IEaOCqZVL+STQ
eXP11L5W8VnodRDh58M/PDksw5YQCFpjJvl8wQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q57uFnCR7T8tBAoMNBT+XJHCC8KWAqe0YCE5G2iK8KpMAdetvYrZDijVNL79FxnPtrl0efDWj6TN
lw/4Cmnm0pJTYWzY4cdb9lpn3rbpFV0yEvHdVl2D6gninJNs0Uz2/E6Ke/cpoUfq2zjpfQ8Tzauw
WBXAcjpYo5Xiq+rsXcmsC1I9ZSkctCHZSKB5JOWh2diBmvO2ag8IncyZ8nMYSWPuYnW8ZlWNL+pC
JE/VTb1mlRKCuy5nI0rEjn+jIPjAhc25VYWaNO9nEipYkzBelLL8JSbsmBFal3yCQaSDwvSBzHbH
4aQFaK/r8V6yR7lJionPar+JhgvyK284MBy9pg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sk2HaHfm82TvnE4/afj3DwTj6+hsiujE5Ltt6Fq/jHWV2t6q59CMzsnceSUKPx4RZIbJl/Q181PQ
ZsmBTBEW9IgLjx5HbJDarOPOz2BSRZIYweKp/8AgCCdYFaAAid2Numa9hGNIMZHX6lEulq5RUE4j
Gb8/nuMc0Uox5TAAfqDaIv7UjUKzaFV/51e2xR3Q6F8Eo4V69ILEHi1N8KepggOJMF00gxvfBbBd
dRKDAPnE1caVZH9Xf42/T+TM0bAwhIfyObwZJSvlYaZceNtLmdudMus9y5jJUZ4Bop4ruUnuGTkx
6q/gbKPwmh//xaA8Hr9rOIz5Ayi+4+nGkX73sw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
p384vz9FHp7DCLW3O/lTGCxfw4G8ZO9oWer4u9Ywwbyzotl2fprbbj//scFDtINQ9aStJOveSBaD
8zx4338oQ5sqUI6+wNoupWc0RFhivVayYKuQ+eKeFDJWQ9eRzBd1iwoZh1/D5/4FzRwFZ52Y6Dx5
/L+yn7KmTMdhpkpwwPw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mvIqzEhj8NgcfeaiFxhx5YejknA/JByLRLxkd2+a+A19X9stdBHzILcp7hfD93GtrbWwYl+rINSv
qZqKWfn4Z4BqupVlmeItUtr61qOV84gMONb4FjVlbygM6fR+jXRLjYGNuQri1Jphak2TPa0MdeXP
YXJy15KUegyU0CTLm3nDHVP0YkPBAAnA2SQ1LHPZmVGYB4RJ1q15+2Awx1zTXPyefMda3Va1wlHz
GdvuKyjrHgEVDz2kSWSZei21SybMnl3IY0ZkgG6ckt+JOtyIl9XEN21FgSMA0vrP8cEwfxPC5PNi
paQ551BLPLze5uwnbrEUELnVtVSrGSD+GTiyjg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 177712)
`protect data_block
ECJVlFcwAZH7B7YXvB8HnAL0ZNFE1AzCMwQYBbF7H+8sqcVP1qHbvC7ABm87je5KFHNJaQBEUTjV
Fu7V6cFPhEBu94yoxBMJm/Xj7BESTkwA1SEavuKWfVIOU/VKCMxV7iuRF8nW/2/yizy9eBPcdTUM
R7ZyugY4DA5jdS2Y1Lu+bPvDOQub3SvEQX1XLgbi+N2RkXB1KSOpHU0f8zXCeZJR2YVw1Plu89MS
Ev+waMjp+YhHjWQ/n9+Ebvg9GnKDpgJ/WivFk5zk+KI4bnvGPoYB3qLNzZ/oiJNpiRT5DPtQcAU2
8bzaQA2GmJ1xxrd7pBZkRXEMmO71G/+E5v9BqZ7L819hYooXRV7GRB+m8eaITHCigfLFfDrLhAoR
2IrkPPt97e8i3PHHpfk5GOgPrb4NK/fFask+YEa5yjzBTQG0v11coQkSTfID/8SzxQZGL2I4AJBT
jHNkOrWBNEuDnWJIdMP/pc5WWld4WdWFRVPtnof9Y1esNXbiHHtAkoZBXS9qwN+H9QAMgqsFnsPR
xBtXRQKXRBr8dYdJP4YkHhIYCX+Z0qjGJCqzHMhMzdFYXdbBD8ChfD66fYHnk6CgSICPaLXsLdM9
bkxRbdt4FaFWZt/OHS/Gjo3EZuOPUXhRXCZUiMAJgius4gu8hwQUxt4vbCKLWrEo2dKiqAXMvAXR
fBrakPn5WA0y5ccBNX8cQPTTf+T7hZ5ysCUGDtnuRj1Y9mDUwXq2E7HE+EYv3VLSi7v9bHaL2d1G
TtUg+gdlxUDtxMXyOdT+GanX9UaKAXWw7J3RbbyJSwxqrTruGVcG7hSVW4eCz6X+swdkNZYvXTur
Rtv5UMDzFYkvxK76b1WBcgqWBFIQU3dDHGGPu0ruJyeh97c13+pSXCqKVyY6llhaQzbzI2k7Ad1p
IFbXbc6izh+0wKk8vfuwcxzfpvZsm9wi001UoEbtlfMU6lyHg6thC/iPvD3apjTCJiHHTO+PjBgP
ZXyQqhJTua9wcek//6btTa0gjrWucRRKtMyKSW2GSpN4/Edyx2he+hQxMf0Ge2RJkMBGuLDmj3Cv
AUO8iOMqqqmMbR3r/vEylOZ4z/olx09uZV6nMeR6xBVLX7l9I6kWSmZtGaHy6hDgeI1QLzIB4m0X
CCMeX7WO3lwtLsjvZOAALV0hEYt+dMJTR0+eQJ5RXzaj5bNFZ7856UZYWfjAvX/tXQA4DTNLEvIF
s2jYhhNU67c9qWgnmtQeWfF5n+nnQmuDupL7Ry1qLraZMhE7nIvXpvTRWbmAMIKtqTy3OXevbMpt
KXsvVmjxfv4k2pVjRpt4ejgFISIGL4u9YUwgR00kqMkdvGkqBFANM/B+bjvMVCQCk+YrZpzsU8s7
ZSL2aO4xldL1TqGQo5rkz/PAHI7HO0mhyoXHtzW20V+T4+UW6YP9qt9gKNfxoofUr70l8w/ImVBq
aFi8s1T1IE6L5XueVvdj1RingWo8swPFXA/c/QkrdOeTi4QU2cOHacUsutxa49qJ9wVVU/0saxzB
685UNS7WvMIV7v/5I45dIxPwIGIE4hVfbzfrX9PLyOl72EOTVPLQBx25/cmUERm4TgqMEyDQ4HzS
wmWodzrvpP2VnZrLoH+NuP0xIn9C2QuyjnIiaL3l6LtXEP6R4M/KmwdwiJaTTb/hNmksu4jiv1cw
Lk1NXTGFsxWG81kK1LWBOtAwSGwpiwzKztLI9WuMgpWVMGEgRSJfCsChCBAYHkPKSNYsTkdpKd81
zCKwd0WLqf4GQaZzgfjCP/oOTS+6WyFxca3DAW+DeH4bJnVN3nK74D0ssrrsoSRbYZU5rc2SpFhN
uHDriO4WQTussyhXofvuqGcJlsJnv2xQmaH27MXV9zI+XF6HVZCDW+9rFzC5SZLtIvQSGmGhtQ7v
6CEtrAaC7jdot0k+T8DKv+cx5uKZ7t1QBLvaRRfSOG6ZIti0VBHyn4lBhxqoWOCdwQvsLbKrzgGf
oqmaOg53dKfrsbVNYAXDgKOlVYw8k4ZkHtyrsz8b6eWAFQ7+0bIogX3aYHDqQM4niZOr5hyO4FgT
0RedOaPIHBiNySOxDStkvlR3sQTnnmHbzQ5Yn2ztXtKKQ5OCZsXFbBHjuE6D8IyKNruRafDFr7+g
eszlphMv6njXdz/O2Jgu2sqAiE29RL/dJGSuos6Ad02ugqigtkEnMDUiE/eFUdwwQ9gpyc1uEiXJ
igRsP7/bq1zDDUrRaFs8LY+o/sj7U7vC5Ku/hOSt7B0xIdsOXgz32Kvf9VSOOELKZezjyhVJ9oxv
cyyQsd7wQTmDPFYs8wKB1kWJhRONqX03w/BtRWvpCotII4OkyJMUY81gQjIYuDieZL9mrl5HLZaK
199VMNHJxDRGzy59REu8dd/Sy/QIdRiRteNauxXWRmV1Avb1IPN6szLOoJJYMtFTJL6TC8kgqt7b
1ni3wII6rcadcWyQCmfgAZ5r9zIR5I7KM+2DTWOeVGceP3H9U/L6A57gz23LCBzwworGVdo2elej
UUiDsK0LDiiwgFTgSR29fYRmvewyCZzKP8ztSoUFmBI4fFsRnJxOyl+X0V7/o1WDZYgYgciMfZkH
rSlhY9+IiMRKKNLhNxMWlHjMCFqSwHqbXkkUZoVu4VXkvnZT13ozvZTXfNKwJVWlp4A4jK9S0USe
yEuQE9JuiLeRnLBz/FdyWx0wLZFjxSQiOoErBjKqS5U38M8+29rntINe/o8ueHJbadFQP2M+fPhG
YHNCTt0JqDshwcAyJjCLMWoAbHJrC5EZddCWZoNHEjX+O12bXeOiJRyDby6W5ZPJ8epEsUBMvTba
CLZj0uqwkJmq1g1AndG3Y2OIkamQywGE/Z1aoeJMQSpoXoTHQFVKIuHJ9xZwzVTG8YObuLwv7A7V
xacBRaH6QyoKREoEWcznso1HI4Seu04V05LndXYF8Bh91kyiYsAywPh6HTarglQHIQaJMkPtWJhY
Oq/4ExunPn/de1YTuf3hFG0EL3tzTs28OXwIowAM6sGAa1IgZ2W6StIUXps1R6L8bIXTGgfi5bWo
yhGW0rsw1vmoYHVM3zV8TqizsHd0guIbTrtG6uO9VJxZvFV55+kFCqe41l4+n73rd8R45Tdx5yi2
a23cigQKYWATXX/OzTL0VLd0Aa2yhJb+SO0WyRkTGchR3aFDQp/HPwclh7fhKFiahz6XeZ9/r42P
PPxKx3mUqQY0zJ87aZFkV41T2z1knCAA2RNyQXhz+OchEhHOFP2XtAdcdTak4oVu4tfHVtIbNGVW
r76obpp/arM/N13WA+aijLXmEqchaexpzRQeocXdgHIqgZnZ8Gna8LnBHF2Ol5yhpy3OIV95Pg74
nwB6oV8CupTjOc9jkoTGF8EVuApKS1/7QmjInaaboQzcLt39TLOsaevO/1Cflw7K5IhA5XkSu/dx
8lMzY6UqAjxhnX4a+heKK1HYjUuWnZg4g6tGgtw3djXl+F7hZYa6psX5WYx9/A8kQZkHpTs5sYhR
hn/AUIaaZ0/88cT5qFEoDqK1d1mNYGMPtLG32cYt6j7eyhQQWEctwQu4StAV0qHdkYWcbu2eKUPb
hBUMgZnu6OWnhT9Y5uhvnBKvmXNfWni51gnugE9u/9AEYp8nNTcy3RmXIBKBNogkF9yE7NjXgbhJ
GbEsJN4RAwi/beW8KlBhIQhXAUOzCKY++UptqaalRIjuwBNZSeQIzKRmDSGIZB2etjRxnJW+r4nQ
dmfghwDzP+MF7M1K5BZ+JJhtKy0bOuId5gyVUWX724ZOepsq+GlS0cZrUbak7ITHXe6uX7oU835J
F6Anb9LrRMw+UNH4CArb+Yv+v4JZhRMg8X/dPIN6NACZ11kLaW3vV8LWkiP5CscMQ2Jhob7PqITS
B1H397qRtJbN9rA/x1UlwDY/z+BYXhUAvBvFG3Eftuinu19RvQUIxKY5t5FC938ZgkiTCXwcKSNx
ebQxKg33Xhk5zMPAVLSxlYdRjxrcvcJY+btyQ/PpZl88r3Vkxg+xcwzwo0vffI0Lxyjelw1GKR9V
E88gWE4TSzcILRJuLXKJb2w/QAPun0CeGIQ7Kft3TWW5dGhygXx1cesNG3kkocFhoQXQdjhr3s8N
mkGRL/Wxun0BWY1vjVy/Fdp3R2Evqq5TpGX6GfmXTAx/lJusevn8oVNf+QPnItYpbJYKvLRBcNTv
fJyfMg5oX6WFk+ZVHQ6+/IqubSaJpRzAATsIiIQM10zjyxrCDeQPACmks6ml8Ez3WqXgMmUodkjx
mQWxpddhc08DNgvZS7MElIsQ9995ClqzmRvh9cmU44c9Mtxxk4BddFtjex7n4Jyo1CaKtd2Hz7kv
0UDU3Gu+LWMDASwfO8VS34FE3SCxR8/Pb69Xy3UPQ71KFVcf1b9tskK08oMBH8fVCYORC61UcZYn
0LERlm76YMVRycKzte3t2tDqNFSJO/cluEP8LYMixE8qhQm85awM0W0jY3L5V2o6Pv9mu2wh8qRr
KiVBx57g+blDmWBI0aVn4Exu8CnrRoKh0BsdoYeP1b1H9TiKszmFJLyvUM5P9jffTGwP2qr7GqhH
6r+dhVZhP21vGmpuZpF9hI2UPQGJ/6CZiMVtDK1f/A7aXaNIwr5m8PRFRrkrxWqFYy8dCAlhl9Kg
Auh4olkdIe1XdRd4at0ElGv5HsLlsVPu0ZwNuI0xxdFZTCxv6JuGW8SukyginvltU6sVX6sD2ZCQ
dtxe7tRYa0adGlW3hM9j/4oWOxeiI/9Tx+tWAmZPJJz4aIZ8tg4Wf9eg/9oQP0mtP3iAw9uC5hiY
qKGyUTr+KbvXpLKehHIqDAJBGvhY9EjO1iyuhXrSe/7e6B2Mm5cuAgY/heNumQAciqdRqvFIEPPv
gjgBKkvR7LozDa7EzDNvMEEd/sX6Y7+M3JlhozUI9uZ4mXucyNAaQnqdGnf5Ge45eXEiUjzuyrOI
o94HvQfGNZouNmzyH5rmq1/FFvRuLpuD1YEhuyfc8IDSpbyWpZKyQ/BOiwY1TEgpZ7eoAMQK5Hm3
pwj3T9kHmOqWcl+PEXMf0naDBrRnVGvyKQKIgBNHkajIpWM8oK8ucvafN8Alm7l0yxUmC0xJHBlt
VWz9e13NdrsJWJKo7x9Q4y3c11WAfxK7cUWbg3FTNsoQ+hO+lNW+6YpO6eI1KJm5hfriEZqBBQ34
jOSsp/HRVOdyfp24c9gs1fSKJzfbv1ceO7icoKppFFDV4QMjsQcQtxx/kPwkofTAf+ftn+p8i/1g
Y8SkcqZpLYxq9ygFWO2g3/jLljPmw5USdPmXczGOriGZe3JCjBlTHLN+NP/7nh2wM/YvYtEGCxXX
Qpc1G7RthI2cWu3NZsmYgH4VUJu3oCMuNv0g9Q6YCH01qtz/HTAfj6zFGJ3LbFATTh5cl61+JddA
gk4sxcK/6S7qd59pv54D9dBy24keYzPfBwqT32ERHr0MG96Q7KPr8Mb+O//te0l2s5HpL4ovkl7q
RrRdke11/maS7pEsjlDhYdbTdsih5l8cQFgz2oSN2AcBeLnM9kK2VaZpwZFLFtsVvIh5n6kFa93w
9mMJOpZGE/E42RcSFRJ53uFCLNebIUy7/JHnWD1vxyJbhSCH6hEu9PWVTl0pcYOPuzUMhkswjO5I
MTNwCF4/XqGKwm6f0f+J4awMOLI8I18rZDlU1biIJWCS3WxAutULObTLe3fKo7LFUtRM34/UOOcn
W8w4dgvw2gmaQiVy26NdSZiScgbw5W0sleIrO7/+bUMI2huhbiuohMk6HZn6oXxfEr6ngCfcrkhW
C6O3qcIN0E4n9TtpxIcmlQBfBHI2wV53pTm4UakoJhfH4yyXI0QBn3UZWNNUWtOh4ZjZ7db2swgB
62t5VvqCqmggpwSdAqHMLVuqgepeo8vmpOlP0MBRHYgam9q4tzLSTrHevFVoSvjad4jsirNEbQXP
7wG6AlQj5WVWlUXxBoVHE3eqEsbv3nOYQ8bwwRKPwMuy+0KvSg2pJ8dHkUcM1lTcvyePHSdYrlor
Qpv7O1eN2rFQN/EKBOAfkI+hZDI7oYmzpjArDxmaeCVirA1RO0yMElC8G/cM+d6u6s8csuzkNxbA
mGkm+YGydRC8GAEISoPzoQozqG9GL736/jLzaodOyVUskgZpdejYEAgivqStIS17FeijyCSEe0z2
Vtls4nT3aX1xKzhdEc9HFW+a2wWEPYdGzMSwhe3DUeF6Na6OOYOJcX4z40apVgfad1yxlkrHY3SP
u8Z+AbKq7kp8Wc5uetEXiQlFKUg1t9d3vrRNRa4+UiHjqUDRVp9BHax5n/9kcrY+KShlyI5MbaZZ
F31q/FCKPOcUvtWRRSjM843yIrW6q4Y5zLwPHYhLS1lXFwj6aq6b6PUwOoBpAIbXuDEyP+LLnzZI
ScMAru0sCN4zV8vPQinLfwgB8kRGcqnur2PnaMUUobcOMNjB4bn4zRkBI+ZOi2eXiLrvlqPZTP4m
h0rK2adQtACD1g9NGb7gpcGKEqT97eHsdunlvOHN6xYLgdT5TT583CYyQuKePLVA+FQm48L83jmq
plfGHs2/9ncYBhy0MTRLTCJ2vSkHtOKFRayGAsSupwcV60tFvYTqxw+szAlbauBFtJ5soDZBMOfU
4tQVIxAfvrCYo0Z3dVl82sqKsKt5xEhka1Ecq8rYujRaJTnfFs1jcX2nAOWHayNlc14hqOJ3Gyld
qbjBvVUd/3TLJo6/wPsyKgdLyDdXMqfq/eBnODgNDpi+X4QWCm+yCjvqG7ZxIK58vnMZBK0WeJDK
Hwi4oGrZItyIzkus+rA4oCBGtGqK5wW3218bTHoiXKb/0G4MavjAieY2FZ8lsDiD7L56E/TPzy+6
QMGRxD4teLMXPchsoXtOXg56mfNp5DYNnzklF43GA13wuyLDtukBQY/crpczOMxd/ROf4rScPDxi
1jRRdiqwOoZRRY0OIxHAGkrGXdUj2Ium5EdtkOZHyS01PpAAfFJkOK2hYAbcTQ+x5CpVDHvByoly
L2NOy4PwvOh1QsM7isnDyke54FZkeNlohbbVICl7KtUkA1TabS20qujBl0ovSRJfSh7GKEgx6JOz
2BRGAHIXWfPdP2rLutJ0qgfTEW3i0+s9pJNNlk6bMlA5nKf5whVXPsePxn/uwIuvqBHj9WdQ9jTJ
/SYA/rp7fWbctCCmCUuL0tnuRmPh7n3FqRFR7dgp45LdD3binZ6ULQvgDs8q9BOyRSlqKU3lGhSf
DJjPkKJ0kZBw6nTOPlp83AP6xquylfXAGtXYHBNmDJjTQg3o2eXarnVWQnZaZNCZ9r7h/AAztl36
XBIIJE9piUb07cAosSJk6z5/Bpsi76xb4pjJs3IbaqXE1Ss+1LXlVOnbUEmYv4AMQoPzf6a+d4tu
lt3hOUCuX5WvNofa6EvFrI06flkPWnkFIJM5pwoiVDNwLH/44l7dqUnZRzeNJTe3uv43Bw/GN7uv
+tpXZW2QjBo7luPwf7NE0WEG+wcfSrVKRQUNo1qP6Vl3I80r8YHWAuRD0DohItEdpVLvM7LSuvYa
RUzmBiwJ2iVF1/bNqboHmxIVV0zmd5hleCBH1dYZl7Vqy5WkiEOXmLnWKE/eU1pGs46XtcC9J6Xp
nEQzdNyUOun0eR6DE5PbN6Q+S0kljihKrN2pC1zDdNkfVaMSYjupHoOt8VuDFH71+js/dK83vxpH
dya64izMYRjMtnYUG/FgxGeHZYFZ22guQe45+8dSNiX2P88u9WXJ6J5c1MEXnjQN3Y2IskO9N3Rn
/fCqrbhS88+R7IptzLXyus5H+LeOspL+4nEHxTusEb5Z12S+jAM61NnEgvRI5YLcNYVl1pdLkvUc
XO7C4GWVuSbhyViZmGcfn5FJ2LcKPO0AnD4wu+gHIRNiz3zvbDX8YiBiThBgRDVeapgm/TaDGMDb
6EZzle8if1HSSUOEuEvhLO7ER1VL1zV2yLVfh69RLyvKdpAX19I3myqbWv/rV+3ye2d9Uu6E9079
hYaGUqPZcvsRKvaQ6wYiMo6xiqfesPa4x7xCrBXMxaBzWeqk0MAesRDOMHk2622ugjFb5CEotpJ7
//6E2/D2cLvG2YepNtwLnXNP6bvbHH13jNmORLzUk/vKUBmo1J6GiIocqwp8zYrNCUtzEZUKBMxj
xXd3oLBbGe0rdDel/5Mkh+62Bd6XozVfrLdKwITqUpQd7t5+rjh3EEEGMV3TiOXdSMdQk7tFdmYI
dHAwdYKd1JO1yMGyNqtW2aVptFbXRuJ/JpPuafooBNGKanGoWE4dp9+ShxxDzdf8ODXWD2gZLS+b
Cbn/ZLAqPWi02/5KOPdIEZ/ADQyFqHx8IYSiE++KQ0rG8asIx2vQJVtpuH+nqKeuEe90FE8hooNV
csGlgUuyhdQXmwi7KiZSga5hTsR/j3R1EZp2jYknufocxgsXy2DB0Rmmcl7mYiC21xz3Rd8XnK/G
5BNVrXpwVzK1mJBKXOnyFn+leJUyKqsvzxCVpzoGf8S5TX/j0cL44H0yDj8Ymkn4D3+5pwAxxvHW
lzCX8q+NCtq4oivzLVpr1jLxEfGZdV/raQSf8BdYEWkW9Jeb69lcwJQ4/x5doU2skSoyvnkliDo2
xrQ6HlLH0YSqyNq+Hf7+alJjX1iqYvU77RSxFfxcwMHegnYJZZpVLFe5xsalnWz5FTvbtZIUh3IA
KZRCREUsrkGHZ9t3+fTUYTLMww2r/1EDnBFiT1ZQtTlfLmi87Bw/rO3EUNhqdRbnkDOENfCBH32C
ksVDLgvIPrMWLhoszIo9TVrpHpM14rodqKz8Sim3N6iDvZCV4cDQds2H9/XRZdnay1R363oMKV7g
p7ACRB7P2/p4d9pip8luNTc2lPD4Q4HU3xTzHVdi/neHaHtQvGOCAtQnY/e+eeqs8/YPHPTAhaBT
cC0MnZXFHJQsxuFhhBUmUDmsbH8Ut26QWaZ9M5qS4uWdsQN5wT0eOtvktYHiZnuxITsMDxTdAbI+
gJz3i0P5MAixbAxaP9SK9hJywYZrTONheOtx8qskYSfCJpsUabIrv7FfEanM+acpL1BxvAtW1SB2
SUyY2TVtDP2PBd/2YQNp1XinYEoTxPE4YcAIzU4cjZ5C8wdnwA4S/lsV05lQ2ZvemYFvhhYR2VJN
vijcilv5rSJ1RgY6z/OaQAngUi9OKAx+70TpkgGY3s0+yn38b6XD97dMV39mGxQWUCjmy3Xmp8bS
T2ksjqLmvCyvJDLOz4BacVG5N+s+xkIhJACKTcgI6Gvd3pqRzp9sH4OynhKLMF2REReu0hz7PmVw
GVUg0VV4G0hwbAh/WUH1+8R4UWDD2W2dYo/zVWtFUE3fa32GpLwN1QX4zoQAuuLva+ynLTw7A337
TtY8bPgFlLaHzH1hw1oo+nBsK5DYFOzNH9774YfnaYTXnvmJUKkUpMONSKxuJ3vSHM5BgUwpKKgg
qkbi3dxyigsiEPw/X8eOPaUZwwkjgjmDvqRyzx/Z6WUtbFb/k1W3WEOYU4T62inlYSCqaE1W1DPQ
NTSxbsuV673s6rbTUkCjXu0sYwwIDhEX+atDGTU3lsHb42mO+24nYW9fMDvDpC6JRPfiZFzflcLN
9AzaGxefSEnww8HWbIO1F791XUcPbyUWU9vZ9mUJzSysgsOauGGXGLOeBXeRqcALhT5E61uQSmSt
7nZ6iV6Sbaep3ORZHIg+y7nw1IGkfJeSnCzrt9eNthpbZsSOlRil5wy0xG68AN9rx6nm36wg/fwy
s+gJfOHyeRHJH+ZqZLCXIcXCAmIPJpBkaVmauDDcqIn6rQkDpS7AELGz1Ic6HC7rRhZp2oCcGtv5
zjzEsw3VloOWXKWNzWwLNFJRDYKD9OQeJU/9qNqqCyfIz4RsWdqNozx1POuZb2Bu7X/vIfPD4S2m
WUyEBEFA7rwTGpmYBsrFMTbfXvmN+CRYnAybHInDky8pCLD5NCFltNSGdHj687k7Zez/j0kuWpgR
XLBl10aN1vauKIjy09FXvAekR564ZKwOY/A575tnVqiR6ouUI99xZlM9K5WVaOZ2PwKggLxFsjoj
g4Nte5KR2EEHcM7xsG70fjJEEyu0qDrYB8K8cXGg1TQFzrGYRJIq7J9gzVBzwUBxjgo43AXFD5V5
DAWlZ7elWV46hCJw/WxTs5QtN8PINmAUu103VGkWTCXvle1/+KZbgTaOlhT+i1hUMFF/hk+1BBH4
PEUm/PHbVTnvPJ+FK1r5POJLrYKWBnhgMkCI4nFeys7QD28gkbnH5Ezsz196MG9HC214eJTSJRWi
hYaswl8napO1k2e/hMNAn0F6hgg6sU1b/4YAReh2SmeUNMHpvOs4zEnwEV4EzrnbH7Bky06xQ0Mn
bk7qTOsfvVkIgn+I3mAzF3kSoM541//fmGuqDbqX4mKWQ5cQxaJleZ722XWVkZXW2Ub4Em/IkO3+
+PVdcSBuj4SkopBMOwkjZqgC3oBUO28JEiYAoz3AeVeYOv8Z2lPkETYQ4CRQmfSdoYbzAKodUVuz
IqKmk5NZaDXf2Z8SO+Y0bg8TerL9L63HxIfWyegLIhjuTpkrEnRYEbKNU5ha0b3bNGipLXfNes0L
7DhSjK4nK81Ky9ep2xGqBNg8EyaX8Tlo6aQaAfZX2b6bRAfZJ5ZJyG5geKr0LG9xNSEotOYrgQHI
N15bq/PcbqPos/uPmkQUqdbc6U2FHmUlLCb9EER8C7gA8Ddpni9r9FlUoZLlTPkSRyNnGkipqfhV
+9lvun4DiWtpTmwvykQkKdVz4Yf4G40NHcrMVa+Rzm6FbSihS2os5uDBY1ceJsGgoinCINnvvngB
tBo1laHU2w6CQd+h0eXH7tPFuk7GubQREsu3UstpRZxwDWkSojhPlQltS6LVzCIC+Egj3Gv2CHpD
Hsvf49LZ8AbiW2+6EYLo2eHPRLQV23UPgliJ09E9eLcLOvIV5xLcHzmxXJ1pBgaBGn7+Srdbx8WR
nEfjr27tuRQxFKj2ijM/ADdXXjwBvTZj2ozCR3I0mQAW264FXaHUfY6h+c1NtcRbc+Ue+mAijOXh
At1BgXDN9eoYk6HgNjJRMAaKe7QzfuzeLaK2fRH1cTt5ALMM1TBBwqxO8bEszX/q1zppmh+f/Qpv
1J3lGturhU0Sz0I5ClTso23ycpW9WehYuaxqdwwq0iyM173zuC1gRCoDGYDIh/QIczGX8Er3mGe5
OQtMMH1uaTB5lzz+CUy/4vxGuAHEUOJzSsNRhOfGtuhy8CzkCMhtlSc/9ZD23t1jRD9BeASdMFxK
sJICQEqaHzh8e71zorAIfaUrXFq6BQxUSi0eg+bnMMRp0oJ7SsAGe1NDhqVomQiJt0r1Rg+VJNQZ
PyuQucdLZwfHZmlzf7xI2PxGdY3B5mEoqK1byD3vmJS/CE2gq7NhYRkQk79YXuQLqxMIhSEiwPp5
9qn4K91PXuXnsXwAaHdG+d0H5PYUgcKtJJGl0c/Wxs9l5KPqBNKoHbu/7dQMqLmLyw5VS8WtdG6y
feB+Tso5DeTEIIWjPBBorm7D9oz+WVVXxsnmnbymKIX61O2qYgF8DrQCaYDiab7SERJjwjmEBgJT
UE96QVD1RkiPuRQKfpjt9Z15JbnKbV9hSG9Z6mCVuHJEFjiNFg1CCcCEuTxPXh6tsF41Q2pYqtT2
6NtinuG25YDczhZv2lTKzg800NkQ5m2F1l4peDiLuSBQfCOjka362yIjlJ7Vt1M5W65qGowGdGlz
fZU7OPWbnVThbWUBheTIWB8wJ0SPC7AjUAC49tQtas+kkjrN07Ve9/WDBetnUwCQIkinEDAlz+j3
8WSANekn/J00TLmW0QK16wlKs7LVWAbyggxBrVGMozd2XWYnzeDeuEDfsSkAy43dG0ifgnHuq9W1
vz6ULDtUmcgGXGTD7kAcV66otmjSt/mvcuh9iLm/JVT+XM3KtP/KnYUchRu9Pe/75dik/NAfma3g
eVvqn1+Hu3G6XLUEr5yTdzzFG6YrlipnFr9eNYHxgnF2nmpTKxND2Pf4PiPrS28b4vR3nro5yvhn
iW8enH6hqfBsDMgety3Hnh4v4qbf9ldGi6LIHDZ0Wzq28WyBpAIE0RmMOhUdxSOtOWu8sfUC4Dp8
jMFuekx4q8OqNMCCIO3edTqcc4GvjT1MEr1iSZMqwLiSK23XOy0ryQjxamOhj8IDbqT1vEN/LEvR
PKasByQxq2+5gNElvqPP4iMZUsz/nkZFdEVFb+lc94BKb8rX07mNe+EHP0n1vv7f+AhNAB0IC0n3
9IhjZIi4CBlZQuym/aPRnO2HoL30V7Lo5FikAmLRe1pQZ2q/V72hUH1Ce0fNp5TB3FfbE/2J4cxo
sW6jdxMTTk7zjBKu6M7Gb87+R6RAInSB56p78FsvjMDqknu0YJ8e5Yt9CQAPQf37thEK7lI4Q117
Q0q7F4V/fIHFn3yRNa8HYGlxcRDVoa46F5vnETojnYbrqPIvNit3gwYYNppzM0+lQVH9/GDpy0Oc
ACZ5TDAI0uBbPuNVQ5zLrH8bhSiQURbwQ4Qu0ep08rA4UawsHcV9LO7iBEnU523WPGex7+0c1ICT
Q0LCd0yOJKuNJhElSmwPKOVu8Kv4iUlcyduUPwcIfXdMl5ay1oMLkSSRm1OscysFwjkeaSOr4kMm
iI0MVSdXLzgAtsN0YIOSdbhxHT5l8MdqIrdYTMm5pZsIbEZn2303rqWWqQ0JKIPN/0Ox/jepmRvC
un7KgMo5uqpSv9Nw0jwfkhczLonUMHkefBqjXKRpTdc9ytkZEWzEHVGWl0t1SsB3Lb4mmeJ06PES
0l1Ml2e+GdO03xDYCLVdCkOmiQD0e5kVwJVa8LhsmiD/iJ9e2OpYglpvB+AmQUzIT5RWgykJX7R1
tPZm6x7fv1zBFB6MCP9mSQ+yUat4832BeoB2+QFY3yMX05bcZEN6bp5cCSyTRvYqOybJ4mw/gbLh
k0QjeHIO5+GAgjvpYOFF82WUoSa8eYdIL/ZojEQHOlqne3DV8L4VbkNHWkCLm8aTy9mxQUYdQ20R
/Ld6V7HXj5r0zd5ewBexS2CXnIDJqA+Y1uaNdcpEed8hmHX3UTMFUq+eFhaGFUXUv2P1qGRDtwna
HzSKIv+hfoYp/mnYnDAQZScy+7KfxMxaxP+p5AGdSp0ZWsELDtsuiYg9/beg+WfHuRYsxTqEOEgO
dyddokpE6BPu9EjUBNRMCv0cSdR+28t2B3WFr27ooJJGCkK+DWfFUSj3qFpge5KKVmZ0AsTKzawW
j5lMEjmssbmuVmENgXVRLAeBAH4XmZYOIvzCnxqQc4Unl/TmthpRp/v3EiYc1CFmUwmb3C3XbHrl
O47IuaABX8DKg9zVFO/ztcT2Nvl9PZnSLuWDt/3UO7zVT8yjIrhVLcfuta5u6NWH1EOFQPkbXF3y
NaGQZ6oGzlUvJcTE7RX6poYqmlQ/EyOyPZMMkpcREFn5T2biBE6jOVHwO3B7vuugEQSESuWgLcFS
eUaz0YP/HTocs5yJBkkPq6LS1fTOmMa9H1vUVyXY84N114r/GnArO4FBAtbsfXXhdYLlkRSLyniX
dmqf06GaxeRC7vzvBbvRYDtyoVaSJNCZVm2aegEUmhbrZalPWt5mwj8CxsyikXwrlodJ6S9vekKa
w0CxB91LSJQbknXdJzJ/o1Dd+jWphLKWOLNimbxeFu8t6yu04szKwfMQjd+eMnh1BZ1eIc74FNrz
WYBzTD+esKjjc4CLh3JfyFqsSTvC4kGiMa4iFU8WpuKp7q6r/i/IRA/4fxA2z1Wrcng9uA+N1ek+
o6LlMk88TRe4srioOBXTCyHZQgEVRf+QVcF+lJYXCTcjz4XS9kUAqOolhuskcBw1zY0RXqviEGI/
AYhOjE6CqzHvlRKo/B9/vV0dml930VcxzRPSeY/NEEtJrFC1NKVfg8JV0gYE6UZf/oQgkBQJO0lQ
8J/PxaFpqar5L+HRZuQ1QjYD6CwzQ4+1QrvsAiyPKz9QVXvPV+CVX8X4d/xu9fG5BwyHIk4cYTUp
P4p5DinyiykqQIlc+UeOPMV2Rhf1RWwGS9Hcq5O+N2rJnUK1KFxMJJdD2I9FRjW9vtWc0nZLr6Ph
iKWsq1yvd/5Ltj64uQm4F/ET8dRN9cTWFdvw/6FVOc8mQLEK+4RTRaUPKFfYoqBQIqDF+s0qUpce
/5/XJpUT1iM3viVtUGqKk/myJT91FC98RMPL6rmBKhU8IsGN1Y7KfLPkWz5IbDcAvHNYyjefFqE0
o25Pj2EBbwou1riiuD7GWXwBfAeZ71d2l4TCA+tWCWD9gvIG5U19nvPCCmf5v4rTIXLP3YA86sO1
8+YQMqMdps5LQRxMA7+5UC3OX6f1gfOdRJEXBl+OfpvPFsHgowicpnIsQ1tkezL6kilaCM0a1X5k
VGsB4NqL47V6+CMLrV1fLqcBJAV0lEVmidzzIbpL5enqOebqRaqU01JXMcSuHMlz4hc3hN/lT2+O
b/ZyqjQDkAxRCg7D07PgPXWYOCrVJWXE/E1DvkuKrvmNajITxrIcyCPyOUEkpzoqpTJEcyY4ZIBd
grZMbiLUUNY1+CL6FfLqQ24Jqvog0wkUdrr3sluCB7kGbBp95GpJ/Fw8w8jWbK4S7DuDHhyn7+Wy
1D4zVG53My3a/QRy1a5EIDpTy7AO2g+UatXpo9P+GZIZfElWljDcJfSO00qf+URB59X8oA05z1eB
cV40+uW+ZK9taLVmKlORk8sNZvogIvz2pupFBEMef9NwBDlWKRM1Dg8CwHLW7UKMEKesuwRx/uic
hPJeHq1frR631fi1vXXL+3+0dkz11m+Ppr5Ty47LucG9qqRZ4lpk5ArKCEcBNC0802ct7y5KsGQG
kXyukK4arx525s6uoojEWEZU7PSN0uVwVQfEk9WZbiOTwnXljHrDoDtVRBpgNVQ/+SZR2MBvevqH
E7M96e7jiinEfXMLs7XHlpEVo0ER0FunhleJ+rZCdxheeweWLQyoSDz+w/v9fkBa+V/G0QgzBhTv
UDD8RpTQtglw6UCQN7aFyegQI+7oC69TN4JFwAeuf4Yl0VdADGIl1vSGvcc5rWYdLl6EEwrECo2a
76QW8b2umU1201bBP360CDMEzsxcJhUGIgQ//yOHjHG8U7bUihJTTe7SF0JnhqyBg58ShY7PDxOy
kz7pz0oS6fNG+HqcOy+Hl8f9GSc5KauGzwM6A3cj7UHyC73ao2U9/65Or/qjjhTm65IwiVmPQazP
9IziDZXVmSUIZQS4eQ0i5+CllLQGPCCRlraMdzNU7Lb1ZD8iQVsFMnT3TrqxJd2PshU5TTryxbaf
rVYKfyYEaZ9PaDrFOC5zJoKb4xc1zNffAuMUGCC//tMhm/acPe+qA3yVPSbs3B1db4DoN41Z5dG9
erhet0lits2z/hc2MAnUqmLFxrMr85eCpcp2YvswswAU19XfwTHH+TR61H12BAUOadXVDy9hf7z8
TnQhWjY2eR3K2CL3PRsuLeHoPnGZBYYgNZTMYuaoYw1XbCMqTTYSX1UVFkgI+fa/SGp3WsrHxj2z
5GNoIhRuSZQFl/0AM0Itgead9ZhPmctbcFLmYYQiiO6mOC+jVbiLXumZclZtdMuM0E7z2kJGoG0T
xBtlMATtE0c+uljXyIxplv9vTQ59ncSaj1NUMzb7wVyXe5hgBPPFfFKnvr28SyqnLC2K6miE+L2B
2wQ/4FypSVMtlp5IxFVNfar9SmXsgVDcOsLsWwezv4xHkYqhZ+PRRVOGbbzBAjcclo7vZhzNfkI1
ynqqH+c06RC5nnAOXxzRchoyAqFnAgbpXrgf1YnFZGrVfg5cl88SJi+fO73ieSasHO+0fRnLkOOd
J5VVAscPoqkT/heziG/D+UE/LpOob4q2gm+i5tjFTGU0rwa1HRjTHKTQ4dZzK+ny2BBkujTIIGFg
UFJw74EEVsnAtMMQ8gIeHzyPUAgXYu6R/CxsWsAxZYkbXezCNe7Quv2P4SOvc005Pvv4f0Ci/BZZ
ccA1DVw9d4I2Tlxm9wVDUwyk9JHyqQsjDKG//KyvkdK0jJvZUHhNE2wmtNpQTxPHw3ggT7AqtgIm
IZ5VufzuWXACxau15bbiURZi57S6a8jse8fv3yUfCcmDKNAsjvY6EhjVWB4wR+3nB1/6K0eMkyHG
MsIJOsoXVF4veK7nptfzO5mgoVgphOUO+Os1/Pj4BYC0nkK2B8YNDfdNMFwCyuHh4pZOw9FpZ9kW
2A+ZbKbgujWVpIA0ZL8PS3QhYDPwxiiNfGQC4rFA1ReO6pRrWt6x/w4ob6YRrFlxMEsIyYPDM4rG
vX+hecREvJJMtup4OTpqOdTp5N35GBCY8akDGcKM4F+grXFfKTDrNt1tZmggM1DicOozKjBYZQCo
eGA5QZXc3Kc/NCoh4d99Zu7Utja0bPobdMQSU+wiNhn8f7NCugYgYIUaJqacbbHt23DO0puEpDgV
qth26B4pGp78ZJKXVF8vpDhS6Fga1t4y4JKI+EyVPO/ygLtyCbK6YY3ujEThUriiVQd6Ky11mpYV
zGyDvgGY3hU4nHuMBuWvqCE1SJfgXloGKlFaeiTqRmLbqgTb8+CqrUKxmi2OyE1LfiPQrMithS1H
wO2PzsxHcDp7oRdeQnr+vSzapUc3qpv6mPonDkMFjExhcV3Qd191D0s/Xa82naYh47y3gYDthPLU
pFJB7r1yp3xBoamtJZwiwr/3ru0LxGgqNld9PDPSW5JQFG6jcz8I1lf+dhNYW+h8wQ9EtkOttfMc
Pw5iXiCcTYyyCGIklcZp1F8Xk0+LNtikF10rq2GyO5YMQ7t0uaNARDHgbBPS5FaQi+cPkO130HtT
7NvEVtnZ4ls9P7wie3xnvf1buLHV8DlF20WX6gOBCrtSB5S+Nfwtf5WR8kzyURE0c594a9SKrVRk
4JcCC+8wbzu5Eqd426ZdVZIP7w/RL40dhCAtym8M4yhItIBETZ5SlxdaVXOfWj/lxyDl6Qnhh6se
lZZkVXoBTRRW6/4SpiyZLBRC2Vi1YO483YFJI6UmmcD3zyAmGWJHenW28pQFyII8e6LiS3r2nAj+
uSQ/Wi9PnF4ajB0Jnnf8MhlnZy2dk7JMcddCRhl1GyXGJHU4PKOlwplLXhe8D0XqiqIHYV4w09w5
RFa7E1WAMIaxM+APG9vv3wRiolz9+4HHEfUekBVUOdkHNg536UN1oh/CL2pjRUqdHRji2pRacB5q
bOKPVT093v86tQxy+zDei3HP5ykUa+ZhvrmV++MQLr5eFlqx0IKmwQMYspsC809BLEglnytLlha2
gxuD/88fI2jI0gMQ0Uaen4zTRIAtbv5Tqo70zngSkB/JHQU69h3Vr/io/rfwCAOLtVk6YDjwxVdE
f+lGPkYjY4Xy2ymEDdG7fmJrHTwUxgkderRTOwGF9RRbIiMbOR7UxgLPl/D39xeLKoWIg/iLvOzP
GrZ7CPmrfRtj3O2iL01SJWMyZ3N5icmU9Ovo6gqK1LQalPjbnAZuiHPTEcFgCozWHZQk/PSqzS+X
foberZ+h8gb5iRH8I6yo598nN68+Qhe8mOKS4LmvFT5ktNSvceTlEEBHILzSqwmWI6PjnvRdb1RH
Uj35KI62rYkry919HdZ8BrQgdgoSOPzlBP9y2QcSVTgRFXMOSznPzNRlQEUrPrxo3ZeFq0zV7YeQ
/rr0IgjITK1Y6c9yP2VhhG4OtiXd6ACdx2utYWkB3NgMGFGVHW6GygEq3PLG2oJ75qHB+XBhB+Zy
Sr7SMxIH2+ygOeR0dxUI6P9gShNGyek7cseL0B1C7sZpuzu9ZTjv28kGxL0OPvP//xeP46ufrpOh
Grf3M14/7qGUKKJcQkhawPwi/i+Upf6mk59ZypX5pErgqrGqhVLYPe6gK4/SYRO+HJzKURr/orNe
fsOUBPbQVjVM7ajqCWIkkj7tRfY5lQ6DneVQL10u9WhGXteLuXaB87yRKCxbXAh4oH/LmKPOn+6B
LRktLSJOfmWEAUJctkBeqsZmBQ7Xkt7ZOwNQrN3ZedP/BZIe58/QDBpOF1O4uVHFttGH3o3mJjUG
Wap9VkCum+ZIy95fP0gfaqhYwnhgdvn4PSh1tTc2KpQbbRweB4a+chas7BCU5vAHjqsDC99zhb8w
xXBUVGzCT6SfI2tnbAd4SRd8jiCD+SKUn8AKgLmJHWmeT1RVT9EuMiijFMHjpzMQNIGN80LHA0SX
hfpFNEPjcnr3dNMsUcA68lSi3SjozrUTPODN4i46WHjuqO0GyBHR9AEf+QX3Pw45bjLictOoFI5V
ZHXwAr+pqLYqQvwKig4b4iBQbWOvb4Ukj/jp82Rn1Mj2M1xtb2pNS/OdLT2tBgw7HHZeGS3JfwOL
3we3AqCQgHNY+hMLrkxQ/43USloSomCNPxbg5ImynGh0qXcBepSGuorcD+0fNZxPwGL0hqOfkpXN
QcRVRZ3M74f9YZHs4py7tquWXkBMYfgrHwyJv1rVGkEKE6GHCOLAjUkBowjYM/llZxF6k2Roli7X
Pwqwt8c4m4M4ABR6+IkQxi64/+WGF4QAbFLxiV5I7PbyLT8SDkyAKAfX/GnQJTIVJO5Q1kFkbmvQ
+4p+CJEsgAQkn2GxYOU4LjiUWI1w09XL992s7XJFdMn/jcFyNPSNpWGS2v60SmVm8pRm0lqpU22W
sQ0qjTMN5l7UdTedYLclt9JGiS3cBRFZG5vUfXfzsyMgYuW3DM6RNezemiaBxeh4E7sOcTR1L7y6
RKCKU1iQLs+OlQZNnsHxOMOWc8Gad1DhuX506eQ4cUFde0l3m0t1ZerTVlf5tw3tXRyR3lUA2PEm
9M6EnJmRZEhxaJmw+PkxtnZiDZITABYD2zzWlDseuP/nOIaXdbE4R6ZrjCLQjct4FnFhgSnB8mLB
zn3KFW3DiOHuEuWAXEQ7mhrt5WSducUvJdGxnkE9o2AEG8PAnhAPKe4pEKfSPKJamk4ciBjwCiNO
403TN1tNxzHiA2JBFZoTKhYZtqiwXT+Rd07YEDZ2ZiJKWfrOX1TDreQXpESFClODKeIOXHNReat2
hz4qLusJB6kh0eRKX/czKRunwCUY17cqVw+cT+6VSEAqoxiJ2ubJnrZk2xmWWlP0EVFYzX6I7E+8
XaMs+IBShSNXOrWn/njEGOu+84E+GVPWgnylpD/1x3v3KjYL+iMuiNSpn5w+4/xbxGAkStTF1a8g
Nzp2HocgIsUPEjDCgVDLtwTephVtvFX0s0+lBSSXG2r2mFsWrWgEG+WPW0fbZ93A6p/4TX2UHf22
4Em/g8DftnjyhvSXQPj3ppinRLRzsw3Olirmn8kapyX7zuo7ARGhumdq1qRezHleebcwlndCP6sH
1XhZjoJ5O0l1kCvWLMaNFqVUxK1TO6Rn3QdKnzI5q48PRSgCd7OVlGTEN7E+ACjW3wSJDWh3ZzaJ
XsNbgT+BfbY4K+NBn5+XyaEX9+FVAYlK+U5f4njeB28orVajJEHbTjnig+vbCWobQgK5awVTTWS+
+mxuA/Prj3/8u2RJL0Didj2zntqkkXpSuTvj+LfOXTlKw/DiqPZYfxI2d9b/WVbZdccZ8sy7Wz4T
Muz+WmSufC9kT3ZvPlNZKcpZaDM8RrBb/eRSxw169T9c/NksPgreLW+ylLmLdp/vCI1nNrgafBsh
MRC5OzHy877m/bIMZlWQQll4dcrtdroUaAuM50CYwTOHWzUmtAfkX2VbGfFOTiNT8g/mI45WZNXN
u5qf7bT+Ng2qrwMQUxR9Qu8lxmWQ8sDi8A5l2xE7V4IVvoxP2DgkeQZ+ltkjvPIigA7iJvYis0os
iyn1Z4eRyEep9LCO/944eStf8mM2X0nZzA2Ghqcyr23+s8jd41nvR663JDsa2AMev2wJffz2VfoL
xmo/1aGi2Jwg8DeEfBZ5PLlb+qwDQxfggdytg/do4Y/GEuPdtIu50moMR88p80unRP6Lqlv3s6Lg
5wgq3SPxFDm0p06AY+Gv3tvfzLqvFS35FH1dlh8LAwklrA/ajssoy/Vae5AAyO7RwBjg1a3ew0Zz
V+10DwNt9xeSW0fOYpvkNzyPu5QAWSYNNkiYJNk4/lI7rqXB68jKhu2vaA9FL81Ouls2Rmd2Swkh
LlWTF4CQXwWygbIZKPd7vPm4Hq5Zqr56rcoiyHbmqT62J2cohqZNfl9Kbxfck6rCiM0iZcMk5b7f
TAjUiSawUO8taQi1aAHSwr2ddYQd4kMqFJfUd2j+BhgBI+FYuIJXuNHIMbrIOAba2ngpHyBHdC8q
l3i3G8IBTfH41sVwNq1nd2m0QmgIW/AGJe7jIKaCxXyXlSsvZly5lj+z1/CKUX7oOZmu8o/fL0ge
lJoa4GZsRFQD3UHZsSchPNVrKOELA0c/duemRqhJxGC4uDBNeyh2FNZhUOmPjfs4VXpEI2dmfGr6
tb5nfo8G/C+uAeiDz1VdCmPX4gqTA+X5nimqlWeQzzJMWd66IR9Y/ap3uzJJZFzSq2BcViUJBxPC
tYFcRW5fBEMrLvrGne82Na1+WTY6tYKZ7kVNwq5ZWEKdRbJqS2HPyHUgAO1IBqD/dQOzj8s+yp9V
4/Rg2GWXyzkCJ2ibRMYH+jQJvIz16JaGl6mjOr1Ai33SbMrtz/9vVw0VsC3O+on+0cxe/hoKm1/3
aA15P4GbSc7JHMLwaPQNqjvApHG3Yv9y1OtrMUKnx1uLSZZPdUc4FZ2aMHan1wiFnmn6cmyiEAQD
e5xXUkZcC/rpFDoxEM83Va5HMXVqQsriQm30PW51hPVEQTu/+XoOvXsltvGi3q1WkgWDyViT+qJ9
cE5QKeNMAzlpya39L/lcLS04TT7T3+aLp/DxhdETC1dIuCpBd8S80i9IocqjYWSNv/2fsfyN0XgT
wkGWyYbwuKi2qFq7N4H/cwfYohFttwOpX9aelQavaUj5HujgA2cKxp1Go0+l/2eFOvtZU4yJ9mUU
Z6mmgoVwswwuGuqonb8foXBO9l2rK1T3DvtNfg486koWUlK+W3ZWLOXRg9C4VvlCH38G1MQra7HE
I9CCFIScpOZwD5fJdJJjXmlUZqibH0a7POrESHLfU670eiYWAVgMjjoVoqgW22n0RWHge7MHtnpJ
o20Xi8kKZ+4EdM9BS71k0T5NsRENc3CnQC/os4UW36ZgZBqX2KCpdf/XcO3bMhm79RmjcVwb85vU
eU0zfCEdFuwiyBaNCILclFM1RT8jXjFaMUlXHBS4LX2N6GM0kMS2z0wFbiX4brUBrPH+9DX3g8uf
YzNf26GAT8+ziwmA0h3oKPEM9NgLD8BuoKfAEbjvUzu0k9mif5pgW+jTGPUsc+AhboOq9kbhLxpb
PVIm5S4nuH7OxJTkTVPstfhz23t2nS1RlM0wSBJ+HCgcCADFk+2SbGk1xz4PgLqlBDJKrljU6LE2
Jv3B6JdAv1vcnMYIeb/UUh/SXtqKKe/hTjNMU82bb5/zGIwrdTEymapsOzqyqYCoRYjaXl70StmI
TtH8koKeio5cHmC3lPdC7kCJr5YG5pL33WeIkFktmwtkNiXvMMmQ/IGIOIdTjs+6fsUW/M/HOvRa
pgYr1kFMfdXX6nYtQ9hZT2Pm3XO/0VKMLE/S/c3eCKz00puv6EP6xy1W0iD2MF+Dz6F7UYyH2EgV
JF6doLstkEzegkoiaOZlhq9O8faOFeceNAFic7AK8GrmmD+iFQpgP74BKkdWEfvOl9ogJ3MPCIcQ
NnPvlEVM7CPi2gHOGNHwgF1EN+DFzm3YEAqy+Hr8/+d1PhYEUiofTRMkv1iT6C48t0tT2Pn6KgIE
THJ388agAsig6WM1S+VqATuX2hbnP3G9/oDv5aKDcEaWFHkwLKNSDyYN9U3Fp1+GfoC8dGf9X70C
6ifBoLThf4sTiZQivIzEe4+d4nWdYO+JqB5KMWMnlyc7mR2MmsobC1lHV/FCajdlgPJCUKT7ZIVV
7by1048ELHbcIBODRWIF44N85yKQ0o1K+/NDbcSlT1Q45P6HyPZzr/BUCy+EuXHnJ138dfkjr4w8
GeYUnI7MxGsktG7EFmVRdTjj4XWjhnSJkxJ2WCrYlRE8sgfjcbOyIVXK5NIgPwEC7v5zRsyL+Hf4
goRCjpdDe55tp8qfR5fHAWoi79tp0KvkkTjFh4HKc/fxRW5RubKFSi7B3SggQ97kWDopPLEyd6r9
8R/TTyYc/o0M1bMuvGwatLb9Rgxb+jNAR0w9knFr+Ij5ViTyJGgSccwdKVl/8/4el0aQfO6nkM0B
2Xhjmgw8Spqra59TIVsE3qrbk+yGPb4lm2vqLdbp7wLYYIQVQHV1ZjlGRFPe9jENbsmM+BPbKDLG
1mu96TWNB92nkIWGZn3UzNLOh4OHQI+kR6hfeTrXWwLUkrJu7lutOjnFwDLkoi2C0Fi8Hjxygz9D
NW9aWQJF7a4dY2EkhW9unn4aYaSpjID+GwHBHs4fFuWwIDfLnvbPUnKFmaff9JpJgyS4kZWsX+Ip
LguxRs/75YiPs9Joy/Nsr/RZxBJj/9+kwAwaaHL8zYmjWZinpogoDnjkM681Y7p+k1ZotjPQ/8wy
ACZIa1bt0IlmdwVfW1uRKvwc/PjdprWZ5Uo0z80frLvEQjE48dJ7ukXccY25KdH2PkEZOb/Z1zNL
SXi8GoHng9IXl0+/LTm1o8eCZxhSTGrLfqrLo3yO91B4MrzMhywwEbJdNSLHrJx1X8heNyaJo8Wx
jkEv4UgaN9WGB/jgjGKe+u7BQEvfRQ6WuYidkq5WvjTokwoAq5+lLFV1FqMLMF3FElOfG7ULyIEF
EFbXN4A3dvBcenamPen4wRQE4OUou2hmekGRgBjQvwuXR568g54vXYZFThDc+kaAgJkmnJKPF5YZ
yUsdEiWpeIgdagjnAQ9qL7SWvZ08JC6J7VNDMH7UFaVJ/eJbHM4CZKcAudkHDONyVIFPS1ebbV0a
Ctn11rsMThft49F8Theg76Q/uNHmLsJJ5uM8tuqfBuBLAGJZS5G5mfcoMyiNPF6i4g1/N13qzP9X
hLAY4cDxrRy6xgi0NoZFr0+nxApX4R66Zyk3GVfiX2y9za172X+eahOQOGHLqLszKoJ4WIdq5RRU
xVgGgDnxObTFoLmTm2KDB7Y51iHI8W3vPx0qxK+XKnGlQ2wj9dDPgtinCyKFck9mCIImnNrfYZzd
ueD2yQKhJJX8+VRREZGRAjEzwQ9bZukvkFQ+M7Ynea0qlazjCuhGHTNAuenOuY1eN6icqaxTcrUf
GkBbnfv5/qQv9ufaSkK42KnYXw1Cr2UT52yO/+tWwH6LRyPQW4X8InMhB4Tsw191JfapQUJv6pHT
ksOA396tfbLUf67JzrG9BP/LUJqTdYfOvTmpsxYcXi8Ioa3PmS8FkJKnl0bZpErN1Qo+I0Ob9YBO
QsJ26lecK9jIfoUBFbxPQjDwKDKTWwH07vaq44XyV4GnA9rD/C8AM5cl9Ai5lrBN0gjvDj3qhile
B/mvzBCX9laUTeZSV+nIKkRFOy0R6gronmDaEP3LfmXF7cLHcB5U+KeaDzxzGtIApUKzNYR/Cw2L
hx36RW2wGB28OUMUOWQqTwHx6xRV39VvJ4kGKyeeGME1KuOmd0T0Z/D561clVRG8e+OP2uUjD5io
iQv681FKrNI9BQDEVVixl6+Ddi0TRIbwoS9/TZQ/W+bMklI3hAr9cTUQFfUzQ5dKKJpRo0iNC+8u
QQMCD3EZoohtw6n9oRZDM4aD7IhNxcNGHB5IWsfeuP75dosJSXPu1uKWr7FIBijv3B9yo+CaCmmn
GKq/od5pcdfNbscMAblCcN27RP+ptzREd8vGNFOV8CAgjQLvVcEO+8sJ99SNiIPEaYFDKGAholG7
Y/aWLlGTWzRMy/ndPGs+Vq++3ZxHBruJG0lzOBMTpPviTxl1anakqlHKt+U+jvFNk3H7WsNXpDl/
cIv9NV30EfjiyCcSRVyEaWJKS1blUCS/C8HWWpvBtW5iCSuVils+0R9T0jOHb9cIElaopOzw5NdA
wuZF6WneANXWIDMazrPsvGAaOyTcAwQlE9IQVW1ascv8fDVeH4fnGIhnYVAmFNHeEMCSzRtKSXAo
ZH1JNOlA79Ox+yZPXSXPaTYCVLd2a8aVxG2ZITZTBrLIFqYDzrdvl019EU1iCiZFOhbS+co6nvEW
sJhiyuSwv0nk1uEsd4p1/3eI4d6kAkWqwaYynQlJAG2SMYP0f2D2Atcl0Db+spDuCwF/iyVh5s9b
APxK9sdwZ9g2IoANU3qoKkRKESdL68Dn+vI0eXvQ8aIdrDvkwOl9u8+T0Frr45Mm7BezQzV/H2IL
G/gzkVyziDdysn73ZROxABx1L2MTBW972G2gK0Ur2Vz+vINRTFxJfJwS32kYaFx9gI9odzuRKRvu
lg+akcoqFiw4+/QKYRFKmxWodQ418vBYMBldsD9fhuBMuBm8g5FdrON6tTfMuJ9Ud+73/FVc/DuV
K+oBGn6KDw7Yy4gph1Q75sKm68kGalTI11YLvnb7DdpYt9XwNPD1TyE72Hu83x8dmXYLYEgF+qus
b4+5nHGNChXRgbpP8MrOB8cOWvvutveBfOLsV6vsuJ646EvSEwxnQVn2Qbymge0AlDsflJ5Xiask
ReBocR1jFkDvv3W8NPYJkH6N7ll0yze1mHbcHR9McY8j4mPZEI8PBWXbBOwRUgc73bJ6KqbL6NPw
+Xs8D7CtgJWcFVvIrPyDXOEvgFHqEvZr55v0ilUIcSpHvNK9jfuUz5FZBg96UHjvWq/Qhye6YrBR
QNZFa3+w+nOe/v00km/UnXMAsozG85zbN18A8WneSnDX1ujZkBdSpZZyS3/Pb6NdvcouQN9VqqHJ
t1F/UOuxVEmGbUN+/LjOZDP/T5t1hbey7eZcWNVwaKhIYS+5hdiu3v2c/E76R9jOrI2i8FeHx4NH
Hji7yfleIoYu66Es7fEn/EIjQ1injRcFmR/yBKrIgUVFFILcIk0+cYfDwwYJZLj+BSvRkt3rEIRX
pggicQFvrOanV/5pKi0SILV/BpzZN7U4GWPo3JQoXBfPU2ULj023xNjy9iEZtPbhnQwCMXx11Gkh
rrdBu5Pffqp2kSu91jqgKkr0TWiLyYzgMMFlkU8v4W2wz217+hkTc+hn/9zgv/zfOtDOlj4EyvDG
+FlGMenjdmak3vPzjUAbxndjerzYKcJcsBF1T0xy1QF7q9jL2PBO0b47IZU1IYnYWrWUkyaso/Jy
2w1Uft+PAaxKdabEhhlqAtW3AIa1cHap3O/aAZ7Eh+BxTsI9yaRPvMlJ62q12R1qZk+TcvAnu4zG
Gdx1Pg8dmvRdORgtOOkdOub0luEE592z+b6Z4gxxqhY3QeJ8GSl7lF+gaVYa/eb/waCmjZlQx55g
lsAM6/lZzOvp0/viRw1sbjsQLBI9TX/3cG4kb+a71Y99l0Yex/Bs4MCx89MyjN0z56Nise6b0cqF
S8iPgreDB5gM0nl4JyXkNVJXHPymu5j9V2dOi7czE2sDCxc9/w7dIP6ghvy1+l4qufzTcY2EIbeF
57MCwAWVLY8ne8Ffi3OuxhZGujkUwf1H4lMUAoXLwkZcKIv4WhJWvGokVk0YN3MO/ot9/yx4Bbwy
djrMSZrC7gj6H/tUI/AveGlT1sLjd06BSSd+SYjXlAIKOY6ZgX8cgumj+RoE8FHYC59XJCPZvUVR
d4yuAWvZbcFeTdEczwnADXg57+t6KYP9RIxd4rwuqOz6GFty0rrEMBnfXX4PsBtVFpeEJ7a+F5B7
VE71DQHjOiZBDd2egqM3zDLUz1Iwxceth1yNjyHV9ecCtaNlPL58817RkYeAwxjokr3T0tln2Znd
SWi0RI0KFGk1zlqwz5zkVYsreXGhrv7Lhkhw6QPxriQ0jAaWCj1epSikmJt2L7kyA8btykqdfcFF
choy1/bcufzmDxJseBUS0H39ZMtaigCuylRCH+QV+KP3goKGMM1YNpcRi/WDhhrqzGb5uwzaJiMe
lN4KtDvHnjSvpZ4hJvDB0MKQrwIHRn+Id8/cZFIEGpaRsueVQYJyjE0OKSeJSTLiRPaL6WIjobxr
dc3Sod1zmuiIEv+4VK5lOwzCz/5OwPuCJ5miaqtOUIPDRv5o7FdAjmL6no5xYtJ3aYKTWRsDPCLS
NxA0snmIkdi2y2QEVdz6ihWp3wYEsWC1NOFlCezZvK3wEET0UX7nLr5a7aPfaJGlfFiHLtP+moSo
ceo12A+BnVoLw6wD/IZAdnVtZOaAI50nNHoq7dvkOxq/XTosXds3URzaYXEgTzBOoiQhnWGnqVQP
2fXQ1vSSXZnMdeeyhdpIT8k4tSAImtRuHdRmAWWYxwU/VeG5e2U0Pjc2rrnGTwiiPJMStrwbU8dK
R5X3CeKybhaiteVal7vD1gdFzH83I7qqubazsfYNfgvUFNyM0aXw561BoyOoY+8dZD8otmJgC5W6
D3VlIwpbFcd/3BgZJ4wcvzFpwEDKDPzASNZXcJPd1ljysHYkitzH7Nq8HHthhfpOWFxqT16ZnZw6
akr5EOCsHnPwK/b/OM+LnU0eLcZGZk7/5ZfdwegsJDFaX+6CZbRv8ew3iG2FBZi2iYyRqLpcp1UZ
TBdi9zBAIwsqOdRciS0S5aTmvA1Tr8ickfmgy4gQAU8MP2LW2AlLy5IaPqnspOCWOwS2u3Jn5i5p
tx9EEHBagvbH28KeOF66uk4oasoVctkfjOXUuxTk3do31VLIzgBmettiXC3AEgGsxK3MJLI5fFHJ
lZKEplCDuyp8KsJqgMAt/M6j+uqjiL1avEHB/wzA0RWlg6uHmia0ZmW9CMB23z4dm//3+/Q98N33
4aMDXkm7rTXYin4D+f1y90MowNp2fDTxJ4mu5D8rHBebseNVJoK3y65LqaPc0XUwIjmcO4oOdHjL
MFagcw1fEpmE8o06qrshuKjAH47RkcaG5ff2sWDrcy8iSTPDsGPkIuhqr4OnjRnJOk3OM1OYodVs
IP1jy29GaBGPMt+oS7RrBTc47fiPmJRsDMtlzpMm/kOpIbdzuSxw2dQMnoRHRhCL9Kp+8lpNYmpl
MlZ1zInzQdJ7dH+0+P3H1nDKHG0h/LP16aMfLH1MkRX9kqj7qPLjaNwbuCJsx4VxFOPdkHJPDd45
QZEEGX5dWHzqdcdoq/R9i9I34lurPdkn+TDS2992nAXpzzN+GnNOHaDooEKx3bXSdQNpSyiytQsO
vu1zvE5tsi5+GPPP5AOx7AxYHGwIZsUL/WwbJilKgX8AWWTm7hcggkX9axpeLQSS+kD/lkZFZdf2
atORJgceBUTfDGPkYFWLNh1JNKRJmZB5fZh7lx3hc0QeVPFt/bo+S5nRoA4MJgstejlB21gi3DAt
SfDQb/Bt1sZ9xgPDkC6o1Vf1bHZnY0Tw1wuA1XzCbOaK1lcSLlb/+BvUZd7N/iQReVikIR7bsbn4
7QS50z+YERIP8MF7fz0qgXEOXJEKcr0OhHF8kLDxEie2Uk6meZijyxaM/JBnKJLmLJIJzx6ZAL71
Rm7boCGqU/hV0WvPGiThTZdRHRp6xKOCoemV81HxZEvJMgAYH9HXHs48wPwMTo4KOf1QxktTdyXt
+mq7RDC9g2QoNJ81ndnuRIogaQ+e8V1dKg9DIwneZFh2d1LhTsA/JPS010I/evoWdONnMxvdZw52
aun+tnzE4HI4//4gMeaTrfcDFHbUaSCESQYlCv0cbhtADzwxV8wDw7JIbfCPg6UOJBTEAVsN9/ZK
AWtlE964kPIe8yecmfU7CYJu/8ItDC8Pvct3lP/IAnSHBH3ii+WTOmHhvIyxjxg3LF5mcUAafi9Y
kzMgAMbPnqSnUhQDaJH93AbXP64lrceaojcwjJep5rn4DvGCpXbSk0DzMefdVEToE6ejDfov9Cxj
lDcsbJYNcoHvhnSEhSTRNFgIfiCtRLcBb9MNTFTsXRGWTmskQppj7qs5Vu620VGI2LEiFykYsqNW
FgZWV1xuPAHNRa4LFpmjIcxVPCvh8cJF7I6FSoB7IXxbYC3jr+xs+fQ3Q3PsTBoYd9GJWA7LMZJB
/YxlLw2dR695l/HI7GUSN8fb4DSQ3B5EGhPlMKCYnqkMu278ytTqBFUupKaUz9Ifzx41EAzdrX86
rQfppH+zDqEfd2v+DmVw+qqCCuetNHUMwG80n9q/kUkxJfO0iBNzkgN3adR4Nwtr26s9biZ585+H
vBexDAa9J+PzVA+wWSYjOkX0CD4wO/wi5OGV3tFdOubmvb5HNeRvHH4JTFSdrCGkpJNxpJfk5Lv7
qqx+4spy+OK2XBSqNFR4PFV7Ke2oYznDzhm5eLtICgsMX2N4z1fQP8mg7+LA684XnjuEUDj7Lxqj
c5psZhEkg/6d0fn9yzkxJnKNsZKMQ0kt5KQWr6TsfxjBh3I3xgM+8282ACz16uxy8xGSnICo7EF/
dUoxeCkCIA8Hg+KeBHMC/K2+YxGn9vlHXD0dDVEABxwpLrXU05oeoB65g6MD9YnhsJLZ6440U2XL
YucjeKCg50dZOk/QPgN3y/KNXKDfHsJvfyXCpJkVON3mq3TaicE91POUbrOx3cwS+VI/Ep2Qrgds
djQqsXzQ0+HyUAm5Jec5weSP6BIntZMK/bVKmTgI0GZf/rIGrmAgxoAXb9hD0hzN1HgYLea9wtJD
pKd4aghVw4fg1/qiJwdhYPq/5UX6DgsQJ29zwR+bSo406ikgteLkgS2exXxHO6uNQSanAvO1cPW5
JsdV31O8VY6RoNumeaS0smSG3+UG7DS4QQcWDiozMH+94tz8lgfmKiZAXHdNFeyLhx1ayr69CxCB
1JeFm/nTcnsINK9E8axeZnbkip9btHO//g0c0dJNPFIPwyrI9QgqCAhwDY+7lhtpfw5TNadfYfku
9Psv05qL0/qSZFxBEUTFPRANkfu2Lw76VXnHos+yO/KROOMHor7bHpbHC6ZD6vvJ62a7mLvTWpLU
+z6z+X0AEseb819qB9yiHTRBWEDxR16upIg7KtVRTOJohIDD/LqEM5aRERQsvxqzqkaz/IEgY+Xj
eQAyddqJUygJAwLhycET4VRVMYgSG/AWIM98/dKIU3C37Kzb0mwZrzQUlfUBdE50tjc2BPjNnQIk
Kg4auSe3SE3M2F27WJH0UgjBUOFveBX/tTW54yGt/bDddDVfuE3r3xQ3oaF77AallIZIJKS9ACxD
a4l813QVNZxTEisu9ptUlXUPJpLlxh/JH7lCpR/luSuJm064B0VphpkqAmwbMPstPEGcq1qiOl6H
scyl7ORW+ovGIuUaCtsmLkf7Uzx0nl5K0AN+QjNAWMe0VG0b373TW1k3C9jT/kWMUDS7dWAou7nO
G5wxgRbX5S4g1nEX66bxZGR8aGx7Nq7wCfO86wzL+ZbAD6j3XzNxhyCxjQ3TPQPSKi2sgO9ya9Bk
nA519814TAda+kEEXg7ukBDRyU0KB3we05dILQX82czLbMhGBDiiOsdVLFjkT8ecat0sUPR+UZIM
paWnwDVL1nkhXpE7K4yUQ6gktmhrATK8j+ncDfSmXooczMdPs+SLtFZGOyozztNgCBoQNcbB8AhR
pjRnIlCZdy6IvZKcbn7sIt3l4/tiPPUkatO2s6QTX/Z29VyRMGDPYPQ8LWATZ8DQk3D90T3RjSS7
bm6ZU5SbQhwDSpFeD0p/6paSH1tiBf6jJrAa3ASWLl8v9vv9oaZtPzYcedwgoXti0IfMfOPlP9J/
1InB8ewtsBvr9E1JVz9PHhPT2Dj30vr3fgDvR3c1oAt+xRerwKroim8tyinFzaADL8VkOBUAu8wB
ZIEPll6dF5BiuvVSEb6UgO/lj8dNdR5QIrzl+uiAgS9UgKDXpIoW2Bg2jFxjwSPeh4EOPJmdkG2l
7h0r9+opN9xS6OrxleMZYSW6bJ0YnSAp98uIfok1KJ7UaEjPdjZNDvpF20gNrPINkaEREKEPMJNx
60LmVOi/mK7G+gZnifKdeKyW7hPUKU+idt8WxuPd7ueMHuTBnVtrx6hhiQYNltkbt+p7oN8Ai5oK
vSFfJBp3vdSmH7PkyK6PFvbewa7kojou24pQW+XdJgGtAb062r/kt0iPfYunZYeb82NOujbBdN1S
n4lOfLVIWRmPnJt99CK/TRKdMTiPEW1yXxTbQ7W2TH2LIDPVtXnXv5AoM0kJLTG1QD0kN2mH5m5n
nix8pRdH9csadSyE13fdUSpHbz0H1PwAjSbMpgyTWOUjkhkZ41mRw5xboCGtqtrlH+DYf67iQJz3
EFVNKVGG9SUuvPumUAc9bGEIKSeCIF7U2q1h4fP/MP16XuY48tKDbTqi9J1M+JuMYzJsr2+AtBuG
eoSQKGducBXhms+KSkl+M0BSDkhC2UnT/rtV6Uha3s2ioBp4dTmfmNxsmgd35Xn4UFdiokPR52Ip
xTbIQFZcfKZD/BtGlqPTAXNq2gLiPmYAgNjnSv6sHHc5P8FTMXrxRnwzwxe1ASszKj55uuLo7QBT
iK5S3YHl/h+cTswdspqIEjvs/4c9L1xb06BNS3/YnzNGBtijjcfB7orKYG0YWmIzWee2jTItfC27
uhZMSQeYpOtOlWhG825S+eMuq5ZUlSDgcOUXqgQdXEnj/EtE1Shwo0OaG1j+KBdjfA3V+hyjc1CT
cp+lvsylbf6b+wuEVbZygHr5Juynp0RWELv8bb4KG4h5H47aibiSVAYwFW2SMZS2+RUnaYGTaFo2
tbGL5PRD1iVU+rgNCHvRuqUIr2vTFLANVL3DIfumDxROZ+kks3H/YzHMSZaFH5+vhohF5sqQsgcv
IYdismPun9DYJ+1OX7NDhp97j27CN+d1U41WVT8JXKaLCT1QXllAg1X4p4p657If43nblIEv70Ix
FeHj2JPxX9b0qmt0JiCWDJDLDXrLCoQFOKcMxlsmQbA5UzEMy7rFvEIjizItKuqohjcPfI6BSJBn
ZI3WS0R3rqnyfiAvxexKxbMhWJ8uTS0YwY37tc7suV0+vhH4TNGkDc+NvYD6zH0i51bOYb/QTc2X
Os8M35jeDGj7CcEKZEaJS6ogBy0QYtU1uGPwH9uVQinceR+uGgZD7Q2dgfxBpUbTpk0+VFY6CpBJ
M79dNAwrf/MlxnBTREAPwnQwXv/sRSqyLu0fXNJ+5WqgyHqoLaTuACZ9e9ygA8Iz0TTERRNwrXGL
lQbPHKo5jA6epSqLxcTnEBhPRIHja+Cy5jUucTCytZbIElvvBRRGlr3OiKeWyT6+5trBgeqH0O+B
rua3aPyzg85VHROwR+LmyevztFINTQ+nh42PZ4h54h+hnQZt7lPR9uTgOtSXN3d7ARvHFbBIdN4G
DZqdd7kQiktG4qbchOEl8g0CFIWAblqowWuvBN7NBB+pN7H9xGNbchHwIrHmYWH0N9ADjnsXn5zW
bFph7LtPoduJwN+Pgh4UcMLnYReHV7FntucKyqlEeEdvR05dv5lfs2xlURjMvytSsGyrKwBlnOht
BFQjim1jgEowF7tL8q/CWGe9YuvV47uQn003FgG4/Oro3ALzP7qJjGUIRfALIMRzzmniYRZF4zBs
Xd6XMsUxc/0KayIMeN90BmtC9ml8Sqn+2VkKbGFSIM6KbTh24Gu+rGbG2hZNEWmUjJFMbOxpB+pE
v9T2D+E860B0ut98PbrV89GygYFWXO+QRdktgAENW3ADkYxnEUvL5hfbbOAfZxjOOsB9yHfADHE/
iiFwR0nvoJ4vdOGdVhfRFUUMSpEYG1kXT3KJPnFVLzYr8q2nxDh18z8u0HwFuve8cdGi0Zye9SkO
hWL0c5xp3xH9Y1CseWhRRiQyE69wrlV9D4iW0440rEo9TTGrLSE2zYp/ZbidI3RA66zGQ5XfnpON
wOSxOpsXRkAMzVna9rRNcjzhn0+AXF+L2UzE9AibKcsAkQHP6r6Zi7H2mpsPoLh4/9pw+uun7hlF
FGBBjXNRlfy1ljzmyrBA3DSbVFxKqDHb2vz4UCKH6XUAywZCRSXJv/kj5UsB4PNdK+K+K7LAIvBD
EECTByksWVw3JxWzf4sRerXV8JfnXCZHkvp1zH2ASSvT2mLdtjFw9tfr0rv3YjLcn7pCZJeCmo8p
ldGfO36uOHONVg8NBW38g5DY3Dg45q/da9qHuI2QY0OC6fcCQo72H5IgRh2+LXdB5JZvWd7f+OyU
3q9/LlyuyhA64qUERZaH/3W2hyQOjaERs7HFuu4taptVBMNo0023CqDhpTU0af8oErJK5FtzvGTE
KkMTbOg/SK6/ss7L0GeKFa0D5xJY5WMIa0FSrh4O2AlNdDxrByFmwlMl0PrucLRvRtOno29ODH8T
HZIB0YNyA8ylb3t9+VIxw3DwonMci8TVsmKdeObM/cPFOBYH332z9DiLNrMQtXQ9LsXAc7gBMATK
6NGR1IooTiQ4ft/segle6+IPdpzFKvWvzXryEpGeVVzyfz5diwFlp9H/ZwcAKKcq2huvG0pNYpv6
TXZ5dLtJz4shdIN/qqr5HsrNhRIb5daLb8WchxFsm0nJMt+xz1yiHB38nVfS6e+RZ3hM2iZdRHCP
ylUygXCG/Z4tIA3FsCaJZjNpM3zXG0tCfpAcjvgUgcs4StJ0+9MBTSP4kvlKsMS9i1SXGNzzNgO9
1FhQwdbyCl9D8MCQPBlpo8pK/7lCXhTO9cqL+kJS86HOsI1bqYF/UqzsHnYrUwi2X1o1xVPjOywY
16c4Uy/3/VcgHIDmr0rdJwL1Cc47dW50CBz4p9WQrl71APT9WF+aSdUTLdENuhW8mUTKla8TiX7h
2kYqnRAju52SaCMVByKO+e0Ade/bmgaIioico9RXs5qVz+kmQeNQIGl355M+HsTsLXt79/SLlmyI
aC3eo/s2HIxj/t6jDukxiGkZO4QFb3DRdf8Q1ZT4Dh/rRgTZI3fJ2Relb+JakLX+mT8ICwcu5uRe
dAIorYItyEmrYsgIeh8iJkOg+Ya+DnjTTtWJRv2N+D2ExmcLbfGkmim2x6MoFNKX3jwA36Xx3Ped
8kXdvVolJvJQSkkjMm2gg7evJ7IKod/7MUJSnEq8MwBjfkbVNfH9jUA09bc72QM8pX+560gIFN3t
OTopZig9zQSQsYzqdLyvHs/Qb5zW1j6rWq4LU0VPSC7/mu7g4LnADqQLpiC128m79Q0Mq+WeQMd0
GQBMtjKm8b6YQrwonhLQG+Zbx76/jIwyWVh1tldUdj7Ogx7HxKrnzTF7WT/5Ty7knGvcMq3ciE95
mfFIIM0CMKVofggVDlcOk4vmd+JayIdpv1HFuJ2I1KTKRXe2xUquSUpsSzfS4RKNVczNNSPcbIuY
S2Yc11i0lS/bL6rbnlfJXhKOrB/uK/BbvLAl+7CR30cDTZ7+A/doZmsvHuO0QGOGOK9v/GFEQ1YN
Fyz2iQ6yvSRJIuTMk7t+jL2+mPeVROIVAoA0sIxplKNBHfKjkv9TmkbXCocfaEKSF3Fw+B+ZBknu
Ngnuc2DHa8xJzHrB2E+nmbs0Hkhp10dG4azOIJbI45GTy+pzBNhIZUCooK0ikda+FKTHqeTgdCHp
YlXjyGnwJy0e1acS9t3v1wCFa6PSaCYjgR1MiInG9vnfrrpAhrlTla12obUiEYLXPk64e1UM1eOE
4iBXBruR5lgWLTEmN+WePht06SXN2uU3qKvsdvM+RmrqIeIQWnyZTqLz/gMh2oKNNiZ6TaFO7k+3
TroGKt0jaJAdWBfCW3dIzpGpprwpsLQpUMU2UdNmgb/JazNSb7ibEc2iICK8CE5C8fBkB1Zcvyb2
Pof+u/Bh22uhLzX5LMQJ8gaiTOQgyTNOAVL9OyFg1GFTuKm+DZHGuno6XVnXzIC9eERgDUVx9jSi
onsO7b8tLVVOOvm8uktb3L37BewSbMj39OnuuHhs5gMv6gx2FarECvG9g/Juxhy6O5ju9CIeg3sA
xOkp+gSeCrplL4RzRTvkTkqaUacdvnUtbAuhF0j3lkBCwEHnPXZ1SSaHgxY+iA7WNCFOpxlud2Pz
6p04OqfAMX82q4UVfl9N4iLQo9+rqVaI3B1xkWABvUml52KtIDlic0MHuKbLWmjJ2AV/nlaZfnwB
Nh0uYH89rihsqPA1hMajHRWT6ACkVecIxZt7AyXSN6jEQ9j4rwcZu7aRPRKt2MoyxS56WqP+KEew
lA+UCJMRr82y3wRLYCJ9mklbLIyiKyXbKr48h9s8UVb/358Epql8lLjX1FFcJIS7cku70bFddnvC
7bS1Tx3wahAy6Iy9+hZ1Jl9gDWRtaYVfVNXOMRuUhZM7/l3LskFVRqocXyv6JMLuQzMrLNKyAuSd
uD9QPxjCiEXbiZPYGBBgiiZ3fHTTC74A22ze1ZbAtVMKe+StZQy1Qdiaew+yLzx2/J4oo6kJpt5+
G6O0nmBGXGk74AY3Z+SEozU3Aibgzij5ZXQxqI4vOo8YaLZ5splkbtMD+uBl58usApaicD032KqS
Dop4pGxUg1MclBgvSldBGN25Mqvobdkd3/cX3h9N6aGlJnAhpww92b/NvGCsv5NEey87i+HC6yKu
Ds0kEG0/8ZEr4Oc8evMxuujid9fCvE1nJ6vQVlVUFikvPIvii0TxtUbjktsUBQ/EvRnQkUGY9Zma
EUtwHKInRQ1A0zzjuPprv8d79LwWK1sg9p/Qv7+DdWOAiLRWWFLdNPr1Hhne2W4CGsIncBScglCN
TrHCpY2mnmFCxPxbzOKq2olLI2zxFg84X0VcUCcY1wUug8HtkLFGwyRk52+1VX0CDKZgn7g8T0qh
53ePk/JaL4qPIa4K+xgCUslMxb/EhkZV9iEwZEb+WcOaEhtO2JrrgTHg5+aFOCFNwAvuFRjVj8eY
vovLYgY0+r3y9f69Z39xGiUf5TE8ig+1NU0VNpZj12ki5VjTHHe8AD9wmVsIdWw8bVEqIkrM1eV6
nmluoOCBp3RBBrwgtXnXjgJxPy0LKceWdrDqDsbukqPrULRZhESDZzXRcyw7JT5QE/1LtQKidAg+
kT/pYB3J3HNcWGaiep0XYUcbyxu29k613vBbIc4lyTcf1oW7qGz8XBkEslGXx6bxk0D/CcdIRhr7
Xx+/0ETf+hwdpn5fL5yVDIqBAiwDXUfN70PCZ3BbRqipmOPqqUSL335HgiVrGLOnEW3e9YI9bjns
3GzzxSpgfod5Pu87M9WC3Ghs8/MUBy/ZFAVm9fAQdqxAW7L8knrhBSckt8Ktqho6iGJ/+ImZtC+W
CpXCR0jHQozL+OSqZKJkBizcl5i6k3KX2uTQbkE+B4DzVOyVTmM6ZmMhMdwD8dm6YdfrGtIcXn0t
WGKN7HzUl+c4zmDzvWYg6xXV08DzMGEo00GfKx5QOZ+vV8XbXIp/9eP4MtN1nC6X5GdYjnQhlwar
Nkt5S1LgYpAgncgbScsCW4ztFeNI9iDIYbDJ+32v+KbqTD/f7/TgcH+qAgnIeDjT9S8JjHVOJM3I
S7Q0ZSw0drAe24cSivqknYLtr9USBBFcblPgR4gnIO1aXnTX56V/v/Pqv3ORGEMWI65jGimY9xZ3
vsHjqIEsiK7Kq/T6uail1S/slIdefaqV9702EPufIqdjWYQhbAivsIZfj4JiaYo5eTv9IDjCJZ3d
hbW+yhTsFSH2uZxwQfaepXDJ3kw2m6Doi821XXAgEQ6HgNBVov/8y0OD8xq3SFRJkY2vMglSt0nz
FgmmIiEvBb/Yp6nOOLu96p6dkcuNBcRXpnfU0IYCpC7vIeFN3gCeKHxDCFaLzjX2kmz6mVVFNlw7
Pge5CdLRw7hivr1rTtZ+w/ICTzeOhjaS+qukihGw0CcaxQCJdaau/3z0ZMAl3IYs1RqgVHXHFJKF
/5O0e6d4IxLNFu8C0quEvnYk31wR0BcjOxSkZ7GuEMkM2UtWOcpdVUGxQ2zo4g9XX0zLZO1R7EtR
EWz8N+w6TtXhVE4FPViPB6irJLKR2+kap8U0bRv9CtwzUTumn9v4hcGbeNG07RquNWrdJDBvWNOu
tOuJfYCs5prg4tmOoadO3OnLJYwfJabiFshs1sXAaOaQnHXtiGdd2auk20qeRR/ENXshsh4mXuJJ
fyUiTWdsw/IlCon/uIP+VIflgr39C9nodVxeAmJPA3Q85Kp/Y/lJVZV/P2Y1c8yacMhI83C1OGOj
6WGwCswNKrjEyFMXH9jbS0QF3Z8cMnUkq43c+HI2Ys3lr/PMByIhJz7LCz+BWtpj/hjLJn/OjwJF
aVcnAuTfM8rfuWr1djO95bW5+A7TQd3qh+Eb4UoPFQiBJ//xk1khJePTzRuZ8ps8Q+gFrAtKwby/
TTV2kGe6UUuV6CHwTTVYomrKCkVJbzd2Vug7wj/swA7pncFPS13GosXPAFoPV6D73kLPc/FSG6Kp
sqHJ7l4FajNghTEe0tRpQ2NsZXHxGS/WOz++Z8o2E/Uiwy2PyKmCiq/pheR58WlnMYSjPQBb8nqP
3drj91DUVR0moXvibh8oAbI+yL0ISK/P9656Hwd3vtxPV/WsAPQjF7gplVQLNSXcn/5eb+7mp6Vo
rJOfxPbBvNcep+tRnGyrOJvGBlLd/0U4OVphofAzlz6PKacf+7TXb1CvdRj2wTHZAhUhNiVRK3ry
2TyqlGHwQDm15up3PoigyIFq7/uJSMkdTTfiqvy7kVvqx7XhuZQVOOZ4h4VVZHlZsrBbrRdjxTRh
VgJYT0UVduo/VR+yzMX9kzViqFue53b4IY42TMo5hnSJr5k3DP1I4f0NG7G4SABOZGRu/tNvpMBR
eq1hQvOJ1mG53TXcZvkbraCK/jxKj6GKWWw7R9iGqCx+73Jl1CDkePd3J7k0mPUb7X4/2o9eF0Es
RZ8exOCrEZIWC8eNzk+5fJLYpLN5eJivVFW3FeoXp0uE2ojWi1Auz1ZK0cF+lUIgUkq/ESzsbM0X
Ige1gkue6tWtrsJVfabkF8oiHtcHsEtHifiS7oiuSRCoVwKas7UbR9Ov/TN5H4H6rmHQNkCN0jeM
dS7Mx8JokA9fv82nMzxGWOpUJ8yRSo3KP4LNP8TPhZLooRUfRETHaNRHss1D6WxcB5IDlBy7llZ0
ACWy+hLkk4incNZA/L3Z208lgjf43Z+/KB79xJ4wko5IOGWPbyXQLCJpEX6AXyB7WbfbdiJqVVuN
bkKdUo/p5no1ijbSh+fSEDHEik+twPHXCOJY5PgSrPIrtgYmkUNCWi5TduUks1/npSNrLcD/f4bh
RSgaqpkfjSLt37fwcJ4R+h7hsuHaRSvEi0lLv9d7nqmECVVyRUrHzFaOG+c2O+4x7Iss9YLzQIAg
c4Mlr+w2LBaN3TX4Gw9Y/jTcFyRFQp318xvPmxxJdWm7/eBouIbqHCCVemiwA9boopvWvqBjctCX
0btT+UG1xQmbSaeEi7NS2mC8benI4aWRHoy0wXpRGgKhWAJaLEB0HlPjQaeTjBDZfXHYFudxdG/x
RVcrs/xPwEhheEWFTFFddG8/mozNdF66p6ZimJZNRk8jgyyF5Bi7rhNmWTl9pjd6IzjUFa7e++Bn
H1s7c27iqdyoaa0GmsQYSm/vXQe2z4oETvyemcpyMUkwX52U1wMsruPheiT9J56dqizLuCNYYpYc
fNhoRj0Z/aVL+jABa80652wPleOlYGDWP3sOqNQL5rZdgacnaPEoAwrrGodmwsoYeExvnOQP/T53
Te5n58ARoBHRMjopFiK3bZb1cWRpfWrEv8nUW6dgm55YBixrITEii3hDMhPovo36j4DAmhE1WNCs
dvVA8ija1vx9djzHQLdkemEt5Vk9r25In2JlzfxXYI2McsyjaMTAIT+uTgZBK/AT52ubQeANAk+Z
h05pa67kCLcXVj9Fh/NdWBpgImjnjClZxTNN/vJ1p+CRQXQdk56tFiacKjaYHrURLZgQ2VZ2eKAf
v0fMW63/GV930TKJYPVZX1zKHLTkx/A5wAESB8ow2mChtj7dslGl4ExPeA5ZrPTQsvJ64opLusM5
0sczBMSo49NRoSjrxv8PY3QedAxaIXt/6WyH1GGCkTn5QC0MMo+TKvsR0MdS5n8BR8s5HNRPrUQR
zNznJVaLoKFoBudonT/1b1JF7SNeMX+DOW7uJaQXgW2jvot5oN+1b5xjp0J1gXyEE0HCq37Ct85u
bQKHwMYOKVMWQb4PX5hfQiY6jN4SOci4C5RcuCwtG/ZZ3H8Nw0QpsODQTThVP0HxZkWJkn88lc50
K6wfkIrZ7Hj06Mth/s55FkPDsluYIZJPB7q7IjuALCP7vbI0ruZAyTZWDbE9U2YITFcVnH19Efzo
6tB47ROlt8KsNpCVx47NOMY5xvvVW7dbWzGtRLAbNmd0K2iNlFaVaE23sbVCmQjbOLMXxPDVnlQN
mFsqtbOvkpIMlg7bNGdkOicF5voxn757LFaUSdl2SLyA1dE7RuF73HSkBrci/6wbCZgGXGHafJWn
T7ZRcwluvQG9ayxzDJ5XXvTZcU9jC9OL2HzFRdie1/yMihMeiMcN2zIRe7/2uWOiU4JOvDMPZt1j
KkJtPEvftaSfxuoXEzr5pMpQ2jL1i7EXjjDKLMl3IGoa92D3evFPvLXIpFR0o4Q+tzo7mYnaYsiW
qGng6174UFzNbrwNcbAXCncoWd2nAed6osONiDGxFpMX0JjLP0Uj00wBCqbGRGtKRorxMKTGGAup
7HWzFBeZUIU0z1KNvAZno8A+E56YOlMm/v+AjfrlO9uVwVv8Yhte3NBeIYsTQJoJxvBAq9IxEkIq
p0pfV5M2lqVRFGQD6O8IL8txPd2S86lnuXLdCc//G0+LB6g7Tm0IDPSgoc/ThriJy0OvEWU29kLY
Ti7xpgBJjF+Jhgcf9TupnbcTKeJqtMs4ijnfjmgfUYPB3eVtWlxecUFTvFEiG3iJxXbBXoUsT61/
GreS+4F4g5D4DfwWW32G1lk7gqr5GuZzU09PsHclN+4qEaZzVqMggUyoQ7pBMR3Q1riRO1D+kANU
DCJ0VoARBFmOWxOYuP2q5pwHtsaRdPkJg4IlVVmprfUgK6fvoUQVInK1AihmW3R0NGv2RkE9pYYX
tQy9bvEbQWG9OFJSLiFUxmh8qp6Zf4UE//HkcYZRJw2G+BnOO66v6gbwzDOlORsZhXOwqKkYVOg7
IwPr7wZwZxvIJia1Hdxd0o8A+CKmJ/aq/l40NCx5Ydohqd8FstYTkclWgFfG2iCtP3nwpBSjwHPD
osxwkBmANbTjEb2n+p4lkvUJHka8zMv9Z1+72td6Y3k4/XTSUZBU3D6Qa8P2jv4B2e6edqkDbmIH
fT6gFD3vwsO51MJRAGC7m9liYhQWZaj+lpO9dkOVK6ZtBleRxu+nvslEjR3rnwP9pCUhmB8Pa1lc
Z49vBc2zpl+NqIjDZSdMlxhzQuigz9MncuIwHy61Ttfe0vnEwPuizQWTs6S5iesjCDmK2x4RSQNF
J1Is82yfLoiVeiDJOWJKCuDfKCOZCEogxh/o0tgXgbCh1+A6V1RbnAiXPrG0x4cYsimhbXcQTa0U
JA739IbUYNDs0fGrQ6fdb8QQEhSkxUFthoena3o/t0W2uvvUuDuVGpEFapaysKDMRHK8dXrkdztR
YAmFnRK4DH1limX14kdQ3lX9Yhaa9C3AgWovxyvUFcQSJEE+ERNrTtC+MqA9vjWeOIKcHFhu8E6o
0C1/dCE9NCwZh4cZDnMejXWDLPIOy1F5T65Mfwq8+ZWGtzRybVtl9+etBkwqiL4IBc6JpGwGIlfF
ddQ7CwGMXSgqDXpvGgLYLb0nRMQ1b1pLPE51/D5heTeqdT11fOFU6811WdQC6TyipnHN0Jo3dcJ7
bTlubt0bdD4t4g+6OfjI3s2Xhg+gpxb2tkDkgYY4pmUqiO4+jDqRa6ztYXIrVHcb+BpZFW2+F6DV
1ybhL4q94itEpLIDpQNL7pmz0E2TsLeLB90HuNmisKXmw9oCGVVf0XRPzRc/TbqmgLFr4ZzgeJ9i
t6qrpDjlUaRNk2QHKdMrSeSShCSbKVkPTRp2bywyEIX9vuzkQLO6DgXd6HMjQ56G1gm820JwFAbW
vvABXtqlwFDnQKfvgaEwXPWHktnMQ9SLBWTOYLY4mGcNoYAgJ4hTJ34jMvITr4tocngCPLAurA7/
E9Pbyua3RQ9azemaUP5Yi09V+g1OPUTgkuSxglhpFHN7Zc9iuIO5JI9favNejwNcK61aSSQydXQp
Dm3th0atdjQrKC6vTPjhnJKLj6+CGAhAKuCAGgBKJUdqi5eZXBV0cO0DVyTN3O61u3g/RzdAWbap
OkmBroQ3Z07hUCNNwdXvnqdVG4UwzSmBnEv8v7nlaqsNqG8Ysidhi5quyA5yO6iBTexmvw9UFmdg
bFCIWNuShTDgxEx/iW92/23SyT7mgm98221hZX9BtmfPEs/vjYelDH006C15k41Hlcs1v5bc1wGs
n+GlP90Bil/HYYaHwI14w8sNv+AEsGgUdcNJCQFMFZViqIz0ApTQ1H6HrcYZLOgznmxgPEVJKT0D
13R9RhZXbP2yfzGgUqA2D/zkbEF2jKprI1COGQI8Ew/KJdd+UUAZ0s6/wB2y041kbWt3ADUBiRuS
iaMIFCJ7EgFb7d/RyIaZuyGcNSImte4EihbfyXL/6rpPzPeRDE52ZK1F5BqfJbFo5JlJRQeSI5+O
5/NGW3X2DYHiIUEFSlOTUkI034+xcGAtL2Kzl6bkF3bsQHHM0GcsBm7JG4JUd1fdpu9I4oFkDhK/
H+DGpfcYVDgVlsBVn/RPlzePIv9l118JjesM+XMOhuKvoTw15ughjhiH+RRLXSzsSBhMYo4uBUvD
MSfzUX/WRvz1kWy2H+uJtpjbjQkws7Qf1t9GPdVe2iyoCXE0IkRdAOh36FPPNHyzAEURYZYnXp97
Md8R2OQZZ888P5nsUgt4aA7GPGN9NuLyzhVKJv3qhgJf9uqRVYGSzVT1/GmKcFjHTY1xAKkBXA62
Gxx3SBwoodkZXo0hDFgfuQiITH2hJr5K5r35hcAPMNDFUVUqDIJsEFC+PTybrFmHf2M4eMoQ2WoV
5B0pCG46e0FLLRVzMd6sEp/RYTNV756lc6oDYWQq1y75DPmFA20Etm72U0DiExCeRBbbyX1+GLnW
wQY06b1ibz+Bl+EVyv7ZENbDUUj5lMS5T5P9Vvz43nNt7ruMXwjRww/8Kv8C2AeckQ7NDm7vRRBM
LrxSMmpuWdi3kIOxax/p5w/DUhhkO7YTSGNPlszmxkb89BCWMw8t/2lhJ04Q8YPtN8zqNWjkn5LM
J1h14g20Pdlbq7WeqE7JhuQ2BzCWvx+o6svYop36TBdkkBnAKFdgGMnnnHRUZhxy/fLwq7N/8HAB
rpzpVcp8d1yHHZGX78gDXyMel4nYfnVt21vxEJPXx0io5SZV7cC+9lSeZsw5gkbL9B0nSa4hM0i/
CQgfD9ZFanWiXkRVe4e2GptoBHSBMLM+zphDQChIkUf2IC6JmWbOc0qzWu5/V1uAsOMvRPljdPFB
UscihxwW+kO3Ik1lwePMQ2wRWNR+qe8cEVZSLNT+nvbhmaBB5e/ghDvRJVeI/EOx/owVMOMXDLw5
TK/B+LSNGaKhm/PjUOoFH8TJ9OEFOXgOSC/F7DJ8fsiDZFBWV50ajtVBkhhcajMITB1ljawEJjFf
Nsn+mWgs2kfFyNaZvdDylbzpbPyXYAUceIYIuwcD7Vu47XKJSlB+3WtoDDb7wlpORy3+ekB1fEDY
GiU79tpwe3n2luz6BVXaesQogf/Cg07W5eDb1Xu1abII6AHUEwKAzEhf2N77lUyGsB6ZKJg+1P/j
HU/nxep/jh9/pstBORqmsSRL9lGrCRBPd3Wb0IqIAUvjybk4kdy5iHRhczWZQ3CoU6IPEq3FllaE
LuKVS2Y20Rk+cH2sFZN0paJe3vQYJJwl6H15SVF1v7VdREvniBR+oLlYaXeLLDt/NV3qqwyL4hf3
mbDeln3r+aAo4ukU67MjWJmjv0zbsAZFZ9gLK5b97mv5+UiNWRQE6i7tS1Z1VnFDq8mw69Bf5Nmt
eh8EBSdR1+UdebMKh/bKNTZG+h+1K90bLm1F3UddBGgk822sAi4X7Z9JT8gVFmQcbpmwT2J9meF3
KUqFKX1lfsgWdiGPMwhBqvn+M4VfBJcmxZV9czeGGjR9U517HEELfbTG5Wql4Xv/E+3TlTkKQOoc
3+x94206kgWyWpXnPJ11hAmmxBaqoA5n39icGF5oesywr1buNiJZ+6112IxIVzBgky9r5YRvU72D
VKNHOVQadY3xn2Lgi8ySlgiiR2GEyBjbddGZTwCcqMtYQBq/FXc7wo1KtmVG4gOFxqgbxEvnptGB
d3tOGkXeHt5eL0qnVxJ5HIP6mLGqddzor5llF6jMeOwbp46clLcX8fGc7E6WQtigR1dyPJoq3JC5
N7RfWI40rLaUwOms3E+QzvtJ11jVCEttS6DqgnWtlpYvLCtzZvecOrRLJm6VzTCTIEQUyoCs1Sla
rqrCi4UfpDHhGIYGOx80+lPRj/tchRCGfwPUFDH/nvo+4MhseWeYsaPqIXhD6rlRfzkw/alp1/GH
G7njTcxJBhUWGCzj9pZOSW6uEIcYMGopXs4KTnss3cJtttiuttbWSZbvI+TJMXJCTLWZHEJIdHoM
6u3M0+SHm1vPcP4E7zDtkZeQSQ9JrNTiEIS2nQu7cjHiP/NamFYD1XlIPRjU5rl8T050MGMPajuc
pC8a9ZPqhvFguDcl+mZFavEZlfltz7Wm6zppHtlHwmxM4oKv8AGB8ZSgMEgYbkjGznNVjFUkmvoV
xbl2qFc4m+5BZIl8OvusTzjS4l6Q5KXJesBMG3FUrKuVakSlc18hQrLXWh0Pee1Q8NLbePIRicOS
o20jqzG56Z12ag5oyxR8d8HTm344HOSVUiToo5YP2JnFfOfE5VNtub4ZlhJ2gKWvhx4VQhHjPELh
jFCj11XEvhz9aMgCdLwA5xSqNDytMKE1vHRJww0SxlXpbClbt0V7NlZ7xrtSIMdUN+6F6H1Br0fu
h4R+HhRtSC/eXd7BCwAtO+bSCDV6iP/L1e8DXvVacaYdFc1UjNjhk7Zs5eiZ2P0syLY3b1PHXc0i
49DIjEdLOTs8ifZA0a0TFmyYOmAvHyMKXWkMnGZU7LuVPkjSO0+zHyLn7dMuq9+MqllTQVaRPMvZ
pDE1Zly5xx282C5WXkyskX2LiUHjXjVyzhiXG9MviWk5mRw5QcD9AeJc6btyf5YVj15Yd3oazwwr
wMOb1lPTsUJzjaXHvTTmPEYh2U1uJviFgEbHWt8+XRkOraRP65u59sIvmzTGq//L2KxyWpNku7ZH
PlGTEZdO/5sa1aGtnpw2cxdVMA4EzcvIW4fh/AZiT7TxyTyL12ATkWPkJQ8HqmjvF0yUHeqsRgYu
6Eqb/UJxHlU0xUmQ5wUWx8IOIuwobPC0aN4fgFolCO8OKnkYfm4DAYs7hlnaz3//5MEzax5cwW7O
odAEMc15BylUEtG/va8160JAOy8FOBfVoacjR2jXFjw+k/eJBeedRbURswDJ34+EUZC0YAYhOQUL
o2SFnJtE7+glin45+2+oWbCmwrsYOu4IbfQjl0NZmS8sA4AWGd7IGq4sgd9YzGRZ5nG74rlOwAgx
ViSCkNO9AVdyYogZnk8PWcB6+kzXVGu+bm9vyKuMGsjXlCsvBGBodhQsiSuetwVsx8S3GC+v8Hom
e7dYjh7dp9xvgTcXiZ5R2PIhOD0/3o6uBVocaFFMKix+oohky1DTnpAdjjAh4hA25o9v0ACQPm5/
IpetkaA3x/mHzxPeeGSCFU65TR7GpIDOrKb5p3TfQws3snR/NgJ0nRHYcg2ZEyLVfNJeKjukMGFV
Dr/MJ7onqgXCIdfO7h9rstkFOTjUzkBgB8yRXmSWjJ4m+4+J2OI2EJCDXRbVrmajAFISWsml/i2y
C2489I0JIRqGzyBuoI1XosvgoNYe6bbKC7ZxXpq53jukF67pVxjC+pPdfLcJ30SB3TE1a+Yw+ok7
s+p7f9xR8LpKaAHtXGqCV/l4srYb7/x31bNnT0VvTqHdLlSA3qUP0RLi39UZdAA+rFQty1tdj6Ld
fDpOGaWrsyu0fdYB+gtmUcFm4Mtr5n80r+Pvebc0TNnyc6BH5smyVW7UJA8mGYMTw3kxRpyEQm+Z
j6Sii5FdBuE3sx7HGxO1hYYx07oSegkVN8SsSD0bH84xY+tSlhSf0Si6im37AtMEviZpwgWR3VWZ
KG8Y/6oKezXjqwQOGdd/YDkOfP6/RVxfZYgEB/yK0Gj1z90sebHf4+jqRzaPWaaBT36RKOncPAuV
gJdleXlXheerN/81jiJ4Y//qx/p4Ygvwm6brf9PVa+FwQ7JnGq0aF715WVX9W6gVrUi+8Skr+Sdy
cer8gHqj1x9TySAnv+azp2ekKvnZR+xFngC0lKml42pnC6o4CTdb3ZMaElws6zW80/9I98J3gT7u
9EHN3LNx27XD2v7HdYU/vYSxLm/CCug/xKVyoaNGg5iXJlL6TRHpQBuL+GF6HMIGLmGEx2J6lvl1
ZoVj5VIM8noKu2tZAfY6vIbXLlcH4ZJsCWXO8JNWMwLZdZL50U6kLtc5JnEgvRF8gMU4LikfAlBj
GtE7zZnfWS2PaiMZin5rdVNMbP+tCUM/oqeUXwonsr2fAx71+8MEnwDXxqYCdvl50OMSLbgdCvJ7
EAzIUzKQgToWXHPKrrTYKo39lNSQSAPBhzYkYNv7GCcBSO0UBQRmcnlGsAwtU6EyiZRfCXplGZ1c
qJ6GDL9ytDsqLX2cHuihRKUmvPyu4gVz8rOXDK0YR16zrOU48CzMuBgWVMexQc+wlzxqlYnNcVFp
b/z4sZ27C5upKB0S8AoalbyTyE+4V39wTPZqrPxA8C4JWPmkCn99A6ZVRBjgtKuFhf7FhnygSq+L
3n7hDuOA4E8Fsw6pECBgGbpGHmclRbnklqH/erBtO2OoyFKFeXRpJv+NeKjQsaTQzfoiug/Bs8xn
rcN8WZrwgXBGTtoBaiSmBtoW8FvN7m/9DYRhTeO8x0jZEODu8EZ6I/yVHcDBj3VKj2YpFAVjCaGr
T0JfT4n7Rw1k9xB2xgAeETvklZegq4lkXusvkP09PGP78khqJQ4Zf22kSqqfr9JFuiwlthmC8wg/
f13SiIQvHTztwRNO4hXGFkkphUuGR8SSFuPbthpPJJV0mi7feuTFBh0+dANmnaSAibvcnVuvnik7
5f+39sMz92jap4+nrABl9THKwI7U5YtMB45Udn5zr9l5R3ozaF2uvHIZ3/02rTpPG38lg025UDFS
s8SLC/K+L0bwftc3xz9enDZR+NxogCIAIK4i+J6nZ2K+a4X/dKceMdO9ycVwzQG0yDqqt7TfRgBH
Y1lu4zv2LNRfDNp9WJtrdyLpE6VmeExS083kccsC0sxbX0873URVxmH5jBsEGttg1bO7lkjddtux
pG9QZwsDA1x7YqD5/KMsCFr/WHJ/xUG19RKkauApsITzuWhPlDp6AHBx7bhmf3yLYx5Vc4lBx+48
3s4jZVMCZBwzNl1AocTELGTS6o6T3fIKBarZGEkepaYwj+T3OWQBHGARF3Zu621aFD+W5YCBWYKs
aPwC3QWFBuONCu0YL1CVpkKz7/CNaS6dJINDmkbgNT3TPEjwfdNT5Yi4DtGsmnOqvbIO5RhFnqQS
c7VkIOkgib0fmwSKBZLGhdqBzrs0X659j8vp/RgPkGgZtjcutu3klwdBIcSM/BNP3T8RYlX5eQkN
gUb6IHFFqpFAyGDuWAy3m3fnE1xaC0lZqUgbgu8FZTJ1+opB+octLPSssmWrU70JnsoTfQAw8848
pRJaV4AGce0OM23rHBKkpNkBleTqldSFbOtTsJ8bvMubbgOn0XZQxf/5COa8cus0t9dF8IPCFpO0
M6Z9lwQCUwWFpgAKn2sb/Xn8F383//7GlAtHBbeNSEPyskHlDmQ19EtoDSr1yk5sXOaSF+dL+MzK
fPjKgB7eEptOp/Du1+vPYMn2aj7eGnT1Vtw/YpMAooYDGxlJqQRqX1fVBLdt79hOkvqjAnGqCKvi
W33NupNVSE2Nt1KVGh8Cnr83xEeytr56Im23jmEBK72lV5nUuCEnCu8JfJLatYmUdR193gFmsds1
5CmXNY1ab3vpEISSNPKgP7VKdExvea4wHH2ChVEgVmtRpJTzgG4+1e6DE0AYVXvnox7m+EvCdnp2
JUIZneRkRU2IH93ThvCuzt5GyRhxhkWsEby0WvD4jrybWYLf2Mi5enSxodVRUvmEWaApaXK1ObGL
3S235KUYh+ZQymXpywOADZ3qqZnfRflXk0IRxzkk+L0MYYJ0tGPew0LcgVL77CV6GKo36dDzJanr
S+7H/phpZM5U++IZqzrudPBu9yY8cWjiEgLgbq1TGmb0D30hCTdLSB66LkTdXfl6nttWikjkFa3c
/4d9vRNZMMVp4QOlJhNBhtN25E6g88chhcMQFpF0xZMuzXJhPldIaS1WcSnTJiT14v8pHVs+ZRCg
tL92MybA+9rEUa/SIPieDJWiwe0F8j/BN5YGPaIrAz16V94zOlrZuCpr5aKrOaNXh5AeaAEIqIt5
/vp98pM9n92WlBmGcWNzuWlEAJLpji4/dY3qvNLqeBmXHIyT2HMRHGvPUa0XI1AChryxJnQFDX8L
NrZ9j7B6FMTUjqfw40ckj4/2++PNzl5J+3gQT+IJIhKp1JJIJ9JJ2kXi2woXcKya/15BJjgewP6s
IIm8H0dN18ypkSWopcA93ah8O3OO0rBLFOwUaxhgUe7/GRnP6U54Jq+SDCcgCJHQOc16u1BTnqQ3
rCFDfk0FtMZWmpuZjsLRMUZIg4Ncclfn8uOKv3SxdCVEJNqk/P20oZWGlLmOa+TN96dzUuPgU1hg
6ipFgBJAaoThNmRjo5unom0b8lRLIJgHmXPvCh5LXRsUs5jetnWxwuqUGtI8mIm+gLgmm0C4YQy3
/27VnTdmrM8tnPmZB5qHmQ+KTCXTLm3jx+SIi/f8r9rn9YTaLXlBOEGa/kI9nFmuzHGKO5nwtFuX
5L8B7lwPCW9Ss36mvNfDQtLU926zoAwgNiYYhe3spoLy7ZNZvvFfCHqxGtEp2UWNObkWeVopnyfQ
tPms5OPL8yQx0ueP7FnfGJEKuHZ0SYI4mqUEEl7BKsjViUQ/mfNUnvI59RRU6Z5Co3Rp+2fPXYk4
zyEfoiH9LykgddnWtGeLPpRx2vBeVv32b7XCv3JjNx3p1B4tWLs8GeyDzG4VQSMh4+m1Ls2IPFd/
+au3nmcDLcPVWDAy8Yn1+JF7n8BH2k/k1y7Xv7QZ8X2/ZQ9MnaII082j2lFj12AjFxS34WRwMmgw
UTClPGog4XjPuIeBLAD4B4QfLC3ld5ObRU7kiooWHXhXuUm5K+3Ta3J2zeY47G5IEfh5+ePpyOMe
b+MeADlynxmqkhqUYG7B5F8Cz7JleTiGQHGuex4naRG1e63V7De1SV5pE/ICU7AKfNhZCuB0gs/R
2dATiMgCPfrgelkZh4oTznPmCLtzkeVNMay0u4i2lnl201fB/7RRREhmC8SZBVzdqn6b9Dy0unHN
Z5YsL2ORoxdZCh0G+EEoYsCX9IO6JXQiVQSngAh9XcCHnf7LtWkcFUq0yAsf0KwyqJ88wwthIfsh
vqdQxxACtfBISzkPVGca5Jv1lKaVXbGqke2nv5jISzVje0jnTtGLmDE8tvOvQI3uCUHxFPHp5c6b
4LZOP9HOcM/fDvlISkg8A5kkOMRpODV5F8tPt1Qbu1ZJP5IDU2VfLf71rzv8TAj6u7hZbkORO8B2
U6LZSTFtyze9PxzLHIZklMvzlGqVu2Ig0TeDGSSMVVZCPzO1Z3pZWYmFqfvdsZLKqy1uUX1wgZvu
E2YmEpMD3LFNvlQLOg1SSkdO+OsGoGdQKaSmM9NdC6unt96h8v+1eR7+wF28i2Z5YRhyTCpufbOj
eE/wwMAOGU2Qrpqti8IDNL+ofxEmRtCT77Rrgf7pP4hmxW3XgX9banmPTu1QD8X+Zm+iNwg4Zfbs
cxVYWHTSra0w/QibKm0ll4EYyjnE6hxAmQAd33Q8Y5pSIfZ9EYyuO5c2qaKl0JJr8RTc9OVPIfny
gtfggzTETF/oBMVQQuE1jf4wzQXVQBcfuk+K9UhfsdEVqZvX6pgiCmw7g0DilAkfV79p2qcMoTne
JAnHbOf9E6IV7M1XcTQc4SRsJMGPumAm5IUHLu/xZvhtRWB8cHQrlzn+zxVuFaQpdd3FOepCbVeR
8Mz7apKi6Im0TMNgCvYGQGr5hnKMV8ALWTMLrEpos1+tiTLn0DU5g6/nRK9lBZ3nfnsGHIEzhNp9
V6V0DXA59MfJuR9UuXV1elfgGjqDrHx9Tlt+iMYKo8xO5Ujuc0jDy6pZKv3RVIjGVPbUXgm7FpMm
Jg9F8tLKZrlwjPvYymeVYks4L6ClEa4enibKFtf+uS7Y0E2ylrJRwbLwqe6f+qnnlS0n2HJvarsq
GqNWjU52wPalgv5ZA1o3mv2jupf6GmZtRfa2am8T4GqkaQQs87Epvat5+39ZMrix3wBFpscLAGtd
L6CGcJ6pqVSyCFaLmyWWYNwnD+TdzFUeopd7NlMq5Vjka8fpDn4bjuAIQ1y6SOpMH0TmAbAXhdlG
pnXpO1U9k0jzboPfrkNAH6N1FRVSGQwQyxJRp1UCXzXPPITTTxT134tHypRPP/do5lWSoCx4SFA/
aI43huE4uKQEN+pbwJsy9dSC90GFRtR+MNsNECOvyT5BtJy2jRPAsOIAT6vxEktIKiwuLdNh5Q3H
OyOm5n3ItGLH8+arbu0DrzqCGLf4qZufMKWp+SbpmfjLHsB+Sul4A/kNmP9MQJdmqheu0dSUoG0l
lSmmCsjITvYKztvakWgYEzOPy7oTVdQFj+BPdO/tY08KpENrS2cKzwspl8ZxFmA0t+FydG0iiiDL
nL+qBf8aiFERCm0NBe9zkSrTd06IZupvP49k1U5lWvrt9C9mVgC/JFkeGSDJdAH3mtQfA6Yqv89u
LD646K2mLGYZ4i0vmIkVcOzV8xUhIxZJ6ajdxHuu8vvtSlP+4MlrLAz8jrchprbAGBraga/CD/xt
FV/Dl53adKwW7utjhyCTvG3CSbki7tygx4WicahL4NqOpHiMHIHIsAanwXYTsJPHN4gtjr14BCXv
Tey/WsuuNEsAj7tUO+Iy3PdCmu5SL4hdmSX4pWwRSZ76QwmN34KZZNLrdX7A31Zjs5x8kcBwGGPL
EjwbR9vJdPMB39GffDoDtg/qo4e9wsKnBrpfkaIPhZDcXUTEzsabe6Yw76+5DypAbBrdJ3RoPzf6
z7IetAtZVYC49a0169P7wuLbcrbKook+fBcKy/VxvLHFzOQbFXBxqdP5QseQf744cgsbQgJ0/dCT
qOQTsaE0To3KaZpJ7Y6hQtK+lh5MO7O3XNJRYzPyMiKFcJnMJthM/2etgl0uwroS4SigCnurDKjZ
wp1RzyYxSArHEvkM/cqpOSlv6GXkh70jCTJ2AUKDZYJxFrlxRSMBi4O599TWfVnvLSfp/OCFCK48
wiq3jbMG7Pc3V2Fr0aXjpEDZuAe2qT/ASwFsaWa/N2Ov0YYU6DelvwikZ0I8nFeR81aqYjzQ1ddx
aBLqPmUObl7nzc8KWmKti85cXtu3FsDMl5xzQax+z2mCJAq1TsyflwmvEFNGf1Wt6LChA2zBdjKc
6FlJKho7f6sjVkYiovPi7jV1tkNVKy8jXGGpMyltxBIFXCtg0FVd63Trh65cPz6AtkumrhGD/FrO
RnHf6WJ39xqcW2HA3bS8MxHZ1xxd77/rt9u7aHeTWkWWqXOE+CLc0hgUW3fWi901TgQfWp+sFFJr
kMLxrc8sTxlqUQHesDJnlcUlDbSvKya0B2lNbVdeXe5UAOjqHxDLUO/HfBIw2g3fFyEUiSX/AVo6
yh0TEMPcDHeUnaJALwwDPsLla4vCtr1zFGKtBzl+kI0S0FThuplMSDptuO2RvDE5inuxH8Bv+FFL
4aoGiONxARTemjleyl/5FUNN95rv5o3evzgYoaOV3KdrseuHRv6l+rHiRCfnoHXmJjGyg7MYBW4N
3j17ETOkswrMHt7Z/b4QjJZPVFmMrnSyOSShJatFEtohGgkMN1c3x9sdHqANjhKHHfQKu94rennl
IeKpaYD4V6fUz7fuAXjVRjMADdrCAFRoSOaJfzT8U4anIjZvnOtVoo1s6LB9dQR9OJum5i82snjV
zHGXV6OeHZBvVGJvqPGqkQNeJvMsxVEvuswADOhu0nJEo7PLGUlNfqffde600J/7i8TEXAM9W30y
t279J+lZKjmjSDiyDQXknNf/x4hmMsFrJ6tB5sJZSBkzlMs89LRomGL6JpJCxC2ZQZQgEgZLELtp
Eq6JTandPPL4Jf15f18VF0Qrr9uM1NDXpHPymByjBz9vyesmhDZAQmN+VfSBkT0q6lARWtZc1Mqr
T6NzE/h9Nj/hlmOz/RTHWspuqS4lVHZThgy5RbtAfklfuW6XR3dTnb2DXvebYMEj96b+9vGKaUN6
7IkKmhlwFCJwH7Kh65ZiUU7RnccTiGSb0cgFzvMHiY3Y266a0U5MxvaNNwb+99VLozUgM6gHGx2R
aJ3EWbawQy+x8Rf5p+zL1O9MnxpfT2Hp3fj+CA7yiHa06aJkQLlbWh7RJLTTKlsyjaKTzBW95cMU
0TPpSLCoQxCh7Bu5uFbQ8jadFF9q2kWueg5VvwZN2GixoAmA6OcxEFrrLKTwkP0OvM/W+wESZ5Yp
jNo8ox06kQPCYUd+0TFGyAT0m6BeXvXSn145j/uVqqSn5pj1wz7cW072sUau2bK8P/u4bd7B+mmF
1Hw1DP+ayCU8EHfAPWBthRbrly5HQpR93Xx1oYYtWDu0qG2DAKtYWxO5UMrTtN/LUUqzO/WNIzqV
DIMdXrViqcIKiHNtaea3wIYLjPPjpUMD8IeC+rThFuxo2zzZ0tU+xw8kThNTgTrWIW6gN1C0JQp2
TAaO4XuC2NOX8qE2Iji59glPlRyxyefvI5licO8UruUz1RgxBiCUgXgdla9rO7xx5dkFf2rOX4Xb
R5nO+gGpK6gXGARJCBHeHKidyAEDntUkpwGS57fCycKapAPZMAXLDGDAemCCoLabIKUnVHSyoE80
An3MGBZOa7a44LFMzZxyaALwKPyUwEW5z99WcB+sD8IMol0YREckmJjRUh50bfebGqC5gmM7lxW9
aC4dFAYj1MunxjgynVBskGR4JjWsg/QghW0nr5TiPIQtFRRrcc2JOIR5wZFpG6wJAug2yRZfWkSN
bqwR196cBo3LvmgBWOVdvQvdy7OAAAg1shYstQeNnsLaGcYIUhA6o15ROU5fhDeYvr2jCAVUIEwf
Ii7Z/t5G+HA+VHx4wcQJHBGe5F+Y9ivg5kYHJuB7RMb8bRVgAK+Ofv3QheT3Jvl/nH6RpOfOePpg
0fPFv3VQFZFx2+TxTPIz0U7Fsx35DDYkHkiJsaIHobUh5/mD29GtHqwzbxy35khKSJBX2Ufp/FHX
gNBNxzJwrh9XUDBpcC3BdpT7AWHakE6iU1D5CnXC2ibKFwNeouLadSW8HLV+cbF6ozuQp+3SXksQ
GVM0KMBu75PiEx942qcELk6DrCNgxq/TX9XJdBw772h2tf9XDqzFlwP+GbkEmnaKPf6db4LfqMzy
0fT9WgNXHrVUXz6nJCwa1A8vIjnMGEMnqHGc1DQ79dLxJrcz3DGJVZ285HSuklCJiMzF7qjkst23
Rz/L4pdOrbgPk/e8y2wTIIs2HGYToATJbZ0lAofQKxL5W0mO11waaE963rOTH0ldpwSwjI8TdyE9
DqHh+r4Db1VerUvGndkbuw3Qz4cNYQQ+94iNOWR66LlsDL95Q6Ib8aNcWfBYdMkgj9i9vJjt70MA
oEFGngZFG/uPZ0zk2rDq0YyjkHz5YYQPW09ISg73tNZDmtQKKpWY+XBttWU7vk80f1rMFFQC+5xz
VpxXbaJKrNA1eSgjAMbC8V6NkPUp5xQaedSiMPSzvUdKPOzq6oyxTvouftHwTw5aHe4V6QuYKpt2
lao6EOsENyohZNKV2cAAS+Txd75MfWreo4NsL0OH9ncCL+9tAHXuGfOGbpR/IRUGxF9S+KHqOfZK
NT+UDtEyfEcY2J0EwZIuowSQTX3UIGxydiLHWBUdgsabriXr6uKTX+UO9b7k9CXmiOx6P/R5MGqB
g+V1oArGzC18xkTzSOx/FLiAiS5jdIhOdzc8nq8pmiMtE2YbLJuGlOQDCHC+Dcc0OkQabFRTVkwM
9e3A2qA7+ogw7qpw/Qu4KZFbQ5N5QZlAlM6FrlKNPj8pfnpAU98C4jOWt9fl4pOAU2GHMY6rSOpx
AzJuWc02OC1lgRKBNZ7VMV2rImD0h6dFgKFzwGK62B/RDMThwoBkvyDJMDmD0GsDnwbmdFIKXKn7
yVQf2Oj3iGstX/Fu0cW9GCCDmga4Q6tGXVs/4CNL3UyckYkcPPD2j5NlEEgrSyV0g5QwIoVD2dbP
OojU1oO4o1DuMUCyrWmoIdWPyBl/MdJyHwOM0M+G3wvzNzWRDWG1GbZ4KlSyra7x68+eZQX2vmbv
UpJq0WsBA18lD7+644G+nXMEMAuWOyUbItDTdtD7p/sk7J/lRULC618PNZrzpVEQCiF8dIRgO3aG
irb6SzAPt+rXnSBmsWt/KOYjraOFAuT8r4ErfoDOmWY8P2DhnWKXnaiISVPdtpu2XeRmRDxCGsW6
WcQOI6Osen7K9vl5SbMqA3MQKGwHFr2BzCyCaljBP0G/XUXusWCMKGANifszLLzBS5LI0lFx2dUm
BKmcXhVxgkEZNCjnYCs5rhwgb6hA9tcgs5dnMnbMGuy1zuFPnFz9zp0kR/ACyFBv+mlRWbEr7dvO
ywKpgpUS9y0lssvaj0vMhir802V1WuVaRAEYs70IRwJd5zFcl7g6r8wwHtfyX+LepnjrhnLI4VRM
mvNDDbGEnGNF6z413E/Fk2jyU3YpmAmJ+sRuqKNyWuAWdeLE7bWQg2u+a0SAEAiqdWDvYq/VdV4K
EstqfG2pwwDXwsYdnMHvc916FGY6GD1A0m4ywAvnWh/IX51zX2f8uF0kj05qcwtfc2Pp6/6XgT3m
i3gs+zfH5Z6CNFqtuK7+7GAQ7vfxCuYGYcclQezYTca1dqPQEBVHDzA9WFGr5oFpO1ztyGgxc7xB
K03Lp6tvTSTF5c04lpiDtWy90xqgt+dRwESkzXqgGsgBEyOp5UeNhkg1cSql6lJ0L24c3N+cfrjj
SfSomwQuGyZX7IUUMyBW3SuOYEzV+Ab5BK1RFZKetvryw/eXuJ9L1/uR6aH8Yvpgv4fApMKms8ES
8i+XURtCZvPTxE8jMMln5f3suxvb9cDUPNPsvRQQv1dtLCqNyq42G2DfHBh9IRehXpc4+CClA5Br
HJZmBaQA99ylc9+69cV4CXmbGbrFHMZLdFtMFZ9Z1ivfC2HDIY2amO7JKAMGU6wYpptxOQYRryik
oYpFSll+thKmp+++UPtJZqcMl7lRe1AFATgi7VQY74ZpLfPiwnsZxMaD2F5Gco+Q+XMeKdkSYCi1
lQ1gvVatsx8b8DVKkGYHOlPGV6salpMQN663fqcrAZiXdTzeU6YOOuxENIpWexwtIsoj05AboLFo
mc9GFVv5+SSrEaptImYsqonbrcsRHabvD3a1IgXzExTzWBUUbc75XAZBAaDTL2Dj0bM2m+KNoWpm
Np+DlGrFvJx9uPajgwDJSjhjKsGskVtBeawo1NULHSCY+ZPLwFNv5cHoGv1cmaB60rBghBSbA8b1
0fGmjgigpj/1BVXc8JRQf2l6LCyduFeHvZ4eo0VQDbLr/XKwTw04oPwbcAvgIBx3PjLLHmTlWX8k
4chU6DzOZ0XZq5e9w9rztWoBAuncEXv87nPCHDJ68gkqVrc7jqgeUUUQ8PG8ezhozdRurnz7mSkr
RG6b4T/DBTnJXF3Fn8CvNHXv01oI9pnyy7VMeFgAtm/xCWL2nRLtzMSAxwyw84m+x+v8YNGhZ0LM
iYRa6iFhAMRVMJJ+ZBuuurZQ2SOrw7eFzGLhqIC8H5MKvtpRq2KgjjNrNBBfF5vNIIjULVbgoTaa
PFvR51FAlUu1UClOyiZ+DdKdfB4U11IcDU43z12Zyx16j66jEZMXMcOb3xoqZc4s5hpTzfM8dGJ2
5prbiCebPALj7DQYfbBR125bQLppzMiFCqKMCzSvh6BD0V7dFAWI56t4kpO6kNwqbmSpgWrft+8s
O0gEu2JWbiThavEO24bvDfT+Zr3Y7xcCu2MMQJxUFVobXqR1Y9/+Egc/5r3h4nfMjeYfZjiBVLdU
2gftINGscBxva6DPkGK5W5/pmSNX7lbOgf0UYQjaIAtqkjBrKpdzvDa2DXOp3Txnfy8fFa88QpP0
cdjQFK9fvb+v6ypV56SnML5EHlizLLPxB1NdRvwvajLA3vhAZqQc6PUtwHh5epOD5IrGzVwpWxVz
E9ubuScHWStjkVz9TNSajCgWIEA8HyqOt/uf9nnzjN2VxYOmh8zAbOVYMOHHGMbaxMqZrYGdQXgz
/f92kXlvf1RVzrhVjfXzQ33YiBWNEzqS4DlZebJ5iAqaLGbeI1kS+D+sux6wUQVVn+32IMkaK1T/
5NNfo/8EB97Wr6qTCBChIEXEqjOlud3EIHdC9nIdHaVrZiKoeVl10yYaFR0XEh76SVgES18lZAq4
hSTGP04pUN29ZlujaB0BGrK1v6lTtCXTV3ueldfJR6kU/wzeIK/DhTnzp2DaskHaTu1dg69ryiqB
AVGinqN1Ic2FZzcLT1hcOb4zYh5G+MZQgweJoBYNvZtHQ2odJg77RS6PvCbEDu9edBdVkohjhyG6
qT+We7AexgGrx+aw1OIBREnmUeLQP4XVHL7CFL0fjjCoTU52gXfocugbtfDUQYASf/EdfF1HHscv
D/WtzyoqCTmDXEMtHKePrTnIxnBePV1DCfFAK9K1iYFHyUer5kU8cUC1nmfGDA+kvsjEEzsgAjok
OoGuqiN9QivkMD44yc/ZDOYGlP/toOFb8/yTWqUxd4HdqTz7T9Wphz2Qe/2kpVpR2hIXKxLRCbK5
iQIMChabd1swI8uCfJqZBGXQdgMirwrxDhIdq0Ampm2XJ6XgqpwfBEcAfkQnhw5mXkSv9Xru0jWb
igMzGeftkmgP1HMglo+37LXF95RxSMQcPbaGhNJbqmv4C8k7s/bVuRrDjUBviymU4X9tsjdXRGKc
FGbA++TdbCmX/i8l97fQmE2Dv85zQlG2l6mbbX6HeBq2kEAB5PlWUBx/Qa72xEW3gIscA8LZahZj
CEVAHe9fALtuWmvXCpeA4WHDnB9ehIKuZCaAK6kY5VnpXI79UPmsAQWHFiWymSrbsCyYBWmSnlbB
FPE7CX2ce5Kj9XnuHKghQZPhiF0ne8e+VXVcf+ZXNLpZ2AC4/xDWE3fBZXBO+Cg8N77TRJpBsFaH
LhF+AHYmHyRaCBRWQAReU5i4xNyp4wpxXKZhtCWMSr8wmGkoidw+EK00dRa5HICj1J2NF8C6wdFi
YzNVtbgyWhFWugVusg1g7fGASkKVQ768c0G1GvFm0ZPPIuhXfnd7DUpkdGmTFBrFL3d07FZWBWsp
WksBipKSvH9vAys3fnmHiHM600TkqFBSvts+p2IWS56u6fxWcQ99UotbSH8QPHL8Zx/wjDaCHFD8
9CtUWiPOsyNHpBtigImTaO2HgNSmgiNe6ASY/XhMHwvYIZpw9o0YHAyEYspnno9q9ZQ+jJOQ0oFb
EAmXE9apAYNKo37gxe2sihayt+6XKpYghgnuaMZLft+Z7KMdJ+jbzI/DsKKYfvDju9Vph/XssntM
vcgUwYLBJtUsyOvVcXAxFOE9BBkawWsiBfh/C8jTdl/5gqn+UkAaUUZezUCXbr3Zakm4dePIJ8ik
GRPVOVTV0hm74wIMnnQSLvahb9HnHQsnlx0dHhpAFdVa7LCh2T1anuJ4bv/rcatFu5SAD6//ZKOp
651lOqI3dTCxKt6QS/Yx6nrLIsKRPVyLz95jqtmQ/ZUJjChqUl6fa1XJamnQDBOu+vW1gyie0c1S
o6g2URM+u6jMITwzdEgHFfYg0WCtbrIG+4q4P7dni+qX5wH63RAdZusOfzx2e5EPDeOsveH81P+e
zacAmVN85zFV0LUMer0kFyAyBjXjyuaYtIwKd8K5csxSMOOIKGZlJXRj6IwDZ4KPVC1QWhrAiRD4
00ZGBC13TCD4XMbjl9wf4hUyNzoyNl/TplcjM8C7iTrBsYq788v1+aXU/Qpx9qToACk6h6KbGfdt
9gQOLxVHZKIJXCssNoyzWuOtA0YeS/n5cO9f9AS8OjC3HDRmbhsPaysvoNGeu+956WVVIbknB41/
oMCCrFRQShnEhKwdJXdQ4h6QgOGC7lQB8rkt1oJpLFqdxN/ZVPYG7HsBbWkDSHcPFoNPVEBJuFPY
AGtfsyDjHFPbfsVXxJyDgbT9ZLB89bZfw0TmO2BTBMz1nBOBf9w0wcdRdinAYGCwCqpyQf1/dTQs
iVGyh6nZpMrYeuIXOXmQVXxqc1wb+SQIrxMYI3mEwq+clEgpPDHcYREkindXsye4vIbxieMy60Vs
4f03U10qjmCAM6+vZnhcbt3+CPwMQNKvJCY4D0STCX7MqTl2qgKJhXqKsCC+Ut+BIlL71PzElAXZ
9M9EiGlPuFRv+X9P2Sz4g8pLbb6F9BM4niJ4gfKx3CrtOIS9BDzYqu+/8WKASXSJ4H7EHfLmLJn+
SDyiu1utkUc1sfDhKRcrerKwL99ZK0Rx1Vybf9/xQK6bvGzbgWjaNspSVzlE8PQsuK7KT2JylgEO
YSsCZQDUAIhxPzYNcZOzKsfQz7/pdTtcmQIvB25jIcKZMRFWEM1B4Rbz9LFwpJlgn/bhBSPGv/mP
CGQ/PFFiu9cBk/1ShHnDxawdFPYKohfbqvgZj3CvSNA32EMHErIBUPB/6Xmj2XN2ceN1vl+40w7Q
CVIVrC+VkRFV2lb5YNEuIZe+sWTZ2KbJK38nOk5Kv6L6nd0sO0dhQ4VmQStx2PZERCiEHXe1UkUw
nSDFHOQXOoR836kp+24BHAAYpmqHSxQZiJKi/DTofj+4u1eiuQyFfOLPQ0kmiE0cR9/otiyUoNF9
RXJ9TlocLnsKkcE5/DU1VzAiC2GwT7o8hs+Zd+b+XEHfgSHNa5oUkDKD8NMoVAwv/MxBFQULQ4/G
1fRvUJ4Bc2OP0tuC0t1SMq2/XA+FSucNfUigfppsKo7ZmE/JVqfqlrXw5JWwKqnPFWv2nx11UJvw
TEMPebaXcXY6EJmuXIPmFC+opEw5IrM4yhJdjSg846rj74K/m9sczkchsy19leyej802ZjTGl0rd
y0texXY4luv1bgbVDiZ7yF5mmpi8riTTA7GYAhXJ2A6mgCzjANgVp3XjxyeVNnK1kffHBNHeET6/
XUV1OnjhrgQyz97rP1ovVHeeFNqKiIWJJk3K8mmO5zU3/ok1hE7cMYW5eidDK+piYRSUdF+SHHe6
sPCcAy9dopJTJuU1V9wmU6MilQxL77u970GZQDFmufMxZNhdTUPH0w86TvkhVitR3pKiBWbVtJRr
ykHIhhOkeRmxywgYOMBz7VFsNoJQZx1i8PzmtkjoyMDDctvHpQZAMVgiVYhLuRTJQ9py064NNQvp
nkshXG5PJCg9PhoSJpEt+4oTSk5HSNlr914VgeYwonW3e6Os+SzLG3SnAwhZcCFp2xIJIKB94Rhq
f1WgeNPfQyn7sTmsAZ2HlaXtMAHEqa6hp7uOuCJPkGb6UR0Zrr6xZ/8K3OjQx30SrNyfho+jVJlp
+EF1tCuBVcV6LQ7NxKjEnJ9HFtVoPUwm71PlR6SF4/8YbigCjgUo2c3j6cHLg6mcjS2RExUjPa09
WVku1VH4Dq/PTOZzRcfPjYSOBmyuutbMfJlRuosMntGJiWgJxoVr1k3DjndkZkqgU7rAELnXf47T
zJE1NngcEBWDP6bCi0mfzaLWhbidzp7qQM0OsDUj9EDf8J8w2AoPZLt8xvMoKnz2qLEpzAgyTUIP
3fJaF2bKIvHlu08edN1wWHbuvlTxJMkIti5225htqwyZ1d2t1y/LVlOmFXr6Q1JKWB6nrUgKTKqG
sKVzXKpTQeDvxNff49Ul89zz7geePTknUgnqgYfPlFEaKd8iFYt0tKHx34UXsN4a2CXsd5iKhTjQ
Ml+b26zuzVkq4WaGcRw+CvazS7FrjgQINb1Y8UEaZe33GGici4tLMmKDkMtXJGbgIUt8a3wBU1DB
Bjj8DKObmeZPv9lYdWjgQDuDE9wx8S9Lnql71J4hTsxwc1E1YBwyM1cuud8+jVTLTQp0D+VXKQw3
ehXLGpy/gE1aVj/Rmd/47U76K+xjPbnagDAtbzZx4R/eJNEw8xImO0Hj1fOKCD1lGPmmZ4JSwuGY
a6/vIviqJ3rDXqud3OO5nLYFNILb4YGnkkizy/y8fafoE553ZNwdSCravs6L2BP9Z9YJVR0xS4Ak
cun+0knoxAifaEB/PH79ZYJy2Y///Fx+QTaISx7JbGp0sMEDzWeZ/GO7n2WIO8r5rf9bVQj8HpX8
VJFnR6cm3Aqn9vw7etbrM2DB6yaSu3O9WC2aOl5go+aGXAzUOgVF1R50061Me+Z0B0oNcAyS9LRf
sXJ2UN+PTh6HhKF0FWV/VmT4aXtyey03E4TYWYN8jsK2xqkPNPZz5xD/Jz6JAPrMFD+4k4kFmFlb
QTihNU7qr6XcbKAv07JbwW/TerUjVXK5uI9ItoUQc3rSNnBIqXOJQ9c+K3wS0faIswqTvDOmkoxE
d7tWmXR/NLyV0U4WvmX8h1lr7yuLCIi4k097iWk34cyOr8Ur0cwv07hJ4F2vEK5HGzi6hYSCWRjE
XJV1TQB3sclI4XLSczTRvFfQ4rMaZsl26Gb/e6Q1od9tCHYFfhtCJOt+j4BPK6GuI02TuU3F/x8H
lCpdH7hsz2j5J0G7F7jMVgFUqlwf4z2kcSfOC4zZK9kqNheFEWDbDBPlMFbheQ9DERIcTpJkTaIH
940tu5rAq71/1RokCPc/ZTA6369X1ISDAtwtptRX5lBDIKRWmT6QfgoWMD361yEW74pI2qb+jnXN
eHIRLecSp/sWRVfg7tTaeAwxtRg7UZkdoF3LIyY3Iza4s7xlGfebYBC1sBrWVVHzjT9s1sVMguc7
3SD06KQXQvpY/f4djVlUV3WyGQGT1NH0CiA0DfEG99DDS9jpLTSOQuOFRDu14DBs0qQc3UrGku1a
D6Mp38ZOYelUkLr2Nhtl68QShQbeTpZOsR3A8VTnvcPYQe7ztNNb0eMoln8T5JnXv7YG93zcLAbq
98SA+NkM18si6lG7MB8mi4bhGPXiUrjOSTnwTay0s7UoUi85S1ZTOie7LQCMtlPowo0MFipbr8QR
muDQnWGRrmMt6VLxdmPw32+KshIemjd7uF+MHlpy6D1bGM7I+XX+d9N3OZZEQxRYUvhpL3hyFWkk
iW7+d9IhXnWcVPTqWpXgTuwWX6SSWfdk3W3DwFvDaZHNLKFlhYFRPwGlD1pBYAfvJUhdDBN8/MXo
0ZDYDCKyvBm9Ry6H/qOYq8tiU/92k5ba78MIzO+NMywwjAi9ynb8Z60QhREzbjsCRHMoyiCGWrRB
FOGBh3G3QtlItaaTn1YVB8Jg9xqNzHFnnmgbo8E4dyL9fa6cEaIWO8Y/++4DyqSzlLyrsr0IIGC2
1FCqbjnSN/DuwvWi1dtGCDxDZJBSGjL0PTNUDfsg/XLgjmz0h6W/q9zZvV8cMj6iVYb6Jj7GEo2P
5ShRCtfXpwAiZYs6QRuqNb+cnsGmGmW+kNThcAKzAaURLl5zUefZIqnShZNFIqV1kuDYuji9ARRe
h7KhnWOZ0B525x31eN4cpS49rnk0/gv/b5/Dk3SQkU5vMYsRgbrjORTC0AaZtwYWb7m90TZENNOh
uIlROpK2KZ8VcmXMbwf+jWj/96U7KfdMwTWGgZ3Q2oe65FjJRMrte6yDIfWFcCkwc1CSs7/e7+FY
HAmyl1CiBCOjC96sBCyHnGj/IQgJn4tl24mx22rNG5XDOIGvOGJ6Vkdb7JMPua+S6g44+NfHDflp
TLzsISyWv5bgExxah2SDuIZ4tBzBB/finHw7ZyeklvL1DSTNNrhFcARaJiLcsY0t/mxYdul4VgOv
V98XZBl18/Z9O8sA3zfALUV3I+ksxT1FezXLLQEcEgXXiKDFJ6dAW8E0mlTrlepiO9bttPfFPlMR
AsnautNCG/LEGv2q7zv/MCRcZbldbqrlLLwCXclyXGWFkMnfO+mhbi5V36nOltjAjyIZ4U011hPU
IWgtU1lvRO1jzTzIzKJnaqBmwt17//VNY8ANdPSODDRTfhHVWnWaBiEO1vq5I54DboY2tt6MbCwo
2uOQ/vQZhMxqFzY9zo79m4b18Jz4LDMV6fGEMEuijOVe85Y7K+7PTY4PXGbbAWjQhHVpLPaG6ZDy
Zg61bRM0kWJ+bJOjp7JBeGN88oYyDOBB7pyqHUDG/Ofbkk7dmSb/4IHGMXcj9UEq2Hdl80tM5ym9
uabLjdWhvwxXjKyQr9zUA8s+Ln8f0SDko2DfBdH++SbuYOTERYL7rkbSreeEvn1RZ9r9KkbX66Gb
rsVyWbg9/etJT35GyY0NUTu61WFykWOgdaM2ltOp8LsWoqa4QsYpJVLfIKhFSB1jcQ2fOPzJhdvN
HA8o6cKfgHpCPPOhO9DlpCanI6VnakY9gFo7kO8eP4iirwDirZ4jWXfOBnzD/6gmBDTa5Sk4juIV
SAnwC5wWLHYzIpcQkCWUeIPs4/cjqwAYNf5/ur5G6N2NSyj5uK5d9NLRz4anRxaDOri80H7KmPXU
1i1sG+xlAeYI+gO5gpM6lLiZ3bGgSjmZ8+skGs3iF3AwZpPtkMcXJEzYt0qxnaLWnTWn7y9TTple
32M+85u7Cfff3A+U4B+LH/wBiJMbCFOw9BchtKQQwviywUSJsQQ+0+pO0VJTsFxSJN2ZE9TTTKmb
WwHmRDy530UFqGLx4zTnObuutNL+fEmCrFU7fWf74c74khxQyO18p8jgcOfVI/RwayP1O/Ming3f
efkoPEJMPmyp6gCwnDuohjf5tlS8ROdOjEDoKGJtuw+Yo60z4+gIyz07C5hWV9PE04OeiH12zUCy
UhOeSnQH0HCbiHysT33BEzi+T/8Q4k93BnEQ96XMJapxTk8WdXrFnOn9ijGOFgcpsmLPW5C35PjF
SWVjqQySPdvMVAj7timfeThIlqMWvzWnqgZRUtpMmP7IZHQ70fsilSmalb/lNYFylhKgHD9ceJbj
1nKwuxshBBfi+UovxQby+MJfh3mnYSlQmXnboG0iejODncC888RFoVuPuAwQgOiHwHnbCgt9NWrz
A0XSxxkNMed/OaV3suimoiw6wsm/Ei2c22L8EDp5G0mEXWuYf+SWEC8bCagoodkRpMx8XPm5Gq7D
+W2hOOH+BRpmLMNxZkZpaFrr5wYZoaAQCsYmsaWS73pIEq5HEAA2kTjAq0NjtIJASoy4vwYOBffI
7el32Ke+Umwti3Vwndepbq88IA48pTMvzS++3eacM15qBGxHLST6/Ho2r7xQ7SnKQLaQQNLnel5d
/lE+MdDL3Nc4KmjUv++14ndUfagTXLqeWZp8Tl1nx1zaFXxsvOZZ4qNVMwuDBEw4BjraTSVxEMYh
veTLhmbIrOOR3m/F//wHlkX3adKq9ZWsesNLglkrbmcUu3H6OM0BdhxiNUWSKDA5AKEcMW23nhXv
/dkKsxa24plfLT5aYnvkKGMvSLRp+uvBh/P7OfCdnqJiQ1j6JMHRxXwm4XH8msxBFg6FlUopBQ9I
vYGWCSmLS44jH0cY/xoTYVaQ+a+oQLcOOOiug/JyEB7kRbGlq7hbltGuKv5b5qjbhsiZR0qQoT76
JfGMBNmXLNgLurpONelv/vTT6onrlejBzknJuggPtZX16OHKyawCokqqUSsQ3JiKdd83QJtlduSx
1erm1A5qk4CTGjSLFNXa2RC4pxyilwMlZog0mniF670BnlKirZ8rqtgx1Ht/5DU6U7U1WxwhhIR7
jDzZvl8GC9RI6tY0toR6FrY0Tst99b3xA9JQYQepbU2TymSdkDfwPYm/t0MgkLqvn+hXEgCi8VEt
0M+aQEC+2Egnhbxb0KiuHsu9vDFOneaIDgYfKU5yec8Ix5EYkN6pfLoU7Qla0AdiSFsUwKp0qKXR
MlpUWHiv2ZKlRdVH5tvA6nsE3a/hpI+zQPRAoYwntzpmUMX64pwrV1BKi2Ed8znAwcS3fCS6O3BD
KyJP5ZU/2o1bd0Gp0PwRvpSlMbmMwnV0elQS238LGuDh/S+iTR5E3KOQ72Xw6lKExPIqYUv+bAB0
HmVulBan7EWjkiYCYiUa1+9kIBobn7AQxhSB5jycy9wi7hiFWeKJjdkxuQ5Y7W5Mcl1E7d5cuH2Q
X8Q8f2XQoycYaLP2IB8aw7gSCY/R/8oIWBA3Ifm9CXTcaRnhDgjLSqr2u93/LVRc32M0APzuK1Vr
dNHuOC8y6RjdBBHeLYs51XKYB6ZF4YEwJZLNSxE5AO3UWb0g23eAHaxe2LhXezLdIC8UjpwkB2Gc
xBHk+BQgQKB8QDgI7OqZYGbSDszC6Sd2m6ywBu4HxzRrXIwhHoGWRV6MhfXPwT6b/tfxT69cJX3z
FuytPBvvBezXbcTks1bbNheJx6xksh+YLnC9HiXi7H5wSYfYmXRHFtyVue+Xdb/E4NieRpkzMR64
zTBoRz3tGy7rG9Od4CUNpm88rZe+LXMGghMg8ZpaD0qRwlgvj4fXzLcmpPt2D16qSZ6x/ZaZYAuv
70W5uRYomLOI2Cjy4ZBRrHcr/8unjKSZcVo67GA944RvDVzmgh/kp5VtSZxay2r9Cv40spvSdoA4
I09ewy5g7FT78NMtDwZvD8KT025w/M0lrXHTtsO/etj0qVSZdCVeTqBPrU8KAjBfXjnRTu7Vhu43
uHWs5UAoAwDwl+wFiPmSRhlM08RW36N8bSexjFFUr1WEY85o5+6DCxamq/uF7eJ/jSJ9RaZvEgFP
Ejr+J4i1b/F6IAIm3DKGXKNPqpLbS49Wj07E06advXvtTT7nwYxlIfb8kI0+NH3UryMKRDplKBY6
gtuW7e05Qox1dKm1gt5yXy1sdHC09S4diL7qc1cKxN7u1xd8g1JnvWeGfrNPQ1OH8bFZoJt2icLN
UwbN01lktvPr2wsdu+ypu1ABGGikJ4Th5MmDQeaxXxtyI8IQZs/biIB+ZRSD90XDGMbJ0PXTjhzD
DOFjl9mietiJxwZxSaL7G0nPrHfC+kq9dUuf4g7DUd75cNH+6G1XmJqbWDd1cI0IXrgl67k5OJK2
NKFaWTk79nBzoDHkuOUdkD84f42wI9u109eZOkvU09Mmjf3oQq+OhQg2wMvflrSN7/Kxjbw01bog
4NaaMflNpcUfyJVgU37iFZLOPNPlsrXXAX3jrk0IvPIfohzWvxCUU78yzeD89ChHq8u50bXperEL
mkdPsefIPOOyybBV6qhpe/fZmlE4nN7uUSfdSM2PeEDfFy8eRosk6N1o6VOKoi2eBwZO3zcG4GQP
fUy2VeIfhR0BLicaLdNhE7ZmZoRNiml4f/9rw/QBAI9nzXO3COHt0PRd+Yi1oHh0t0MSaSMmvEDw
pTnmPHThsn6jwl/41YKwzhLXeFXqcfKXfUk6LamiqE+uiqPsG/CLbriXri2gUApNxMJqzPOfMxE0
IdXMcF8KXc/5IGw5ONKwehIzGpLgiiQTMe+4XNK5HV54Tf5up+6tVhrav4tzVo737LV0R1KN2LbA
pOVwWc7iP3G8rousVZywujTv4Vi3owWWf8hDaxj763F/57Dw6uyIzcyOW0+rDkExbQtlmFI9dRP2
hwQwl8Ia+0Il4xNEQVsI9KGI+MQhtVuvzkqObrWBJokOXJmNRhRwjK3YhFlqu25XLOoMduHWlWUM
TCW7cS0e4mudQSpLs/GsFAbKPBfBLGzIItsDZvDJC75V08UU4d4MwogCWGvjLkjv8UsEVHMR4RQP
LS567Ux+5s9eFiX90/ANAJhtj+1Y9l/9B7+LGGJT+KmvyFUT2ZQGk+UMdsfa38IYZPXbqR2CR0vH
krMFhev+Qs66gu+rkuA8ymFrb8phJ2LfubRJj4dmcQCo2wHK3xID9l1DhYNaBkBuR1Hbz2LI82c9
a+tqahcf4HIR7KAgb4w2WFJ/6Iqi8jhuJBjZqLOeDr5GtAQQFo5On6vpmN1GPsSdVJdTu0Nge+/o
Ze/zpG7BOF78EUfrzNACiS1cx8Ocsjy8E8/UKcPEA6c9C52ohcvF6UcGC2XOlZWdw+n4Lr8RMzF7
Vtglm9nctNeygGqf9WizJBm5++IMfPh0WHxj/r87GQLkfJIYqu8uGyyD5g3AetIlJSOylcBdyVNH
C4XWJmE8J85r9YZEtAMMgYv2Dt2XRWYOcLVwX5zgNwlIrKYdSYo9qj9aB4jr14pqn3ewhwNYiw7c
Qr1ev5JVuPQ4AX61JKTqTNRa/gfte8XZMC7syg/73nmXBh/NFNZrPmSSsMBGJthhH1//vpH8PHBZ
P222NnQOv3ftTUDMyePyiz0bdCdZ810p5n8cj9Id2I1u7q57KPowfILDd0/w6eeeaN4kEnpZWJS+
CwZTHqMqr55uOIO0bKd1a8NP7ObX8Lr2PWffwwPhTJgrNkaVYTuaIh9EiqEVsNRdOr9+vChJGQqT
hC18yd5czT151nHSYJx+OiplAWFOBO2W8V2fGHHqPh0FxRm5wNay0NuYG300waI1GsA0hcWfqNDR
9DsJbku2nF/+Z9P6If6/+53rfxUEq6D593q5TcKUziwfW2fiQ03wjnLj4LcRFTjbt48k7zrlTfML
bxlM+34qJnkOYkdajXqBc81xqbYwdu9zl0Hrh1/tZDIld97TnvBEcr+CltLhXf9xle7sLu2HWZUw
0A+8sSkGouD2EQrEdX4gBlS7x4HUB16j5n7dF5KThJF7jssEmLMyinqjffJr7cgotcFDVyjLf541
RkY0/ujM0WsiP436HKwFdVYnM52r54D0/E0lGPxpmCDDpfJ7yuOnFHbHSDngo+SUuxV2XXvHax0m
ewiXUVzaI0360IzKZvdx9nQiIImlQJYpW2pobFQjSHozAw9TT+WftDiyLKwAfitGzSO5QZXKA/4C
VTJlCEx6pUdrijs+BBdbIEBHorMDFLo9HQVJhVAFjOrKzUBdKQ25wifxgWSMGUsjgiZUjZIDTfKO
iLtnrNsai/OQmBK0BoE+l1es1r/H3KZkMoa8GA1Ck0y2DxKN9b9QSx8XXOUMYFVoNTh2ClummiXh
oK7C4IBe98cz3C4LR+tiA6LrIh2dWulDRFBqfTPSF9nDX6Uewi9Ve4eqUHh+CQ/sdJtelXIU0Iwn
hEVyjC4iiIlnUboKD/VI1HiuFUKh5f/DvLnl+43mkp+6pnaopfRSRJgsSf3lN6hPoL7oGg05NL16
IcaX/eNqe3Q5niNwGTweu/j6WqCR60si8gxewknzGdLrzwnJ3+AeTRI8AXQozSGadgbvZpQGp5+p
kxcSrcXcr6xr8QXUoXb0IftP0Vbz5k2rUGLXtWv+gyuJ9yFkp6kBl6fwAHofVGYy3lWzQcxrFxfz
L0kpDPZD5sB+wzV+OQVc5AKW4CpGtAYbiCxrh2muQdiwFc69+T3lWjF/aFIfYbocdL6cTT20wTUZ
0+z6+iENOLc2KhTWCdP9nJ747PR2CEE64oDfjMkQFb8slJCgCvMZmK0+tUUXbSaEj0j/awWPdo6I
xr/lTN9bJXhyUb8sVNiTq60/y/L9e/M6n6m8Q3bkopVro+U3RLla945a7ryaJAAWSiZF0OdGEGtl
X3HwtsxRhTuSP55PivYe5zVAJXgPk7cSbgTsz0B7+UicLbchi4DCx2rAzkcCc79pL319/clsDU/B
DFErE+qs71HC2nTUN10Wu9U/Y012nKUXYfzxUefl0tVOza4AeJURdZoz4xEsmlpm9Y4a2pk5EPf8
WPQpfwQOl1WRZffwfEdEcD3u5IPc0YJJk8FBXs5BCPGKVvuj20RmnZpDNjTUJKnUGvTj5tiQBWER
Vaxgptil00/+akwoqByZJvTUSG5h1NTdbSG3pHlucXtMLECkx/KrO/Ovqfdtq0OqYj7RITgSGwuV
XXi4UlVxuH6Q3gOZXpNMCOgos+d8Uodgjwh0sjBHN02LD7WWGubx522k+du1zwveIdqCOBEtFyHH
96PlknRMZIAoz/x4qliut9/A5+jXrXfkSF4pi6auTLX0Wj0yTd4/G5J6jk9hObtU5g52+kJXq04p
ncM/MsXWj8jfO/L165fGkgmSuvqoBXix8lD4brFaJKJpXGJwHoQdbrKWv7dH8vRzq4ejnt7L3sTy
LPupRjNLnVmMXgBipcR2IVHGajvXb6rh71YV6kme8RMG0i+ZtfQBxFTv1cgxs34UE3nhYXWUFCKD
CLnFwKwJgeMo48IMbXE1TLiW293ek1oG9nNbg7/vo3ClcgycaPwCd5wPUiMXRfBHqHcOZKHtRa1Q
8t9lO3lFuVyUCthVbLC4MJarMMOfbNnJud3vJNS3bX0dBCkJF497F8jEViMd25RUFZN5tb+syd4C
fkyRQmEq6q1LWYCKen9zr8BTd09ciEekuZISpyx7OL0+ct10aIRjaJj0kY0jP83xpyL0flTt9tY8
h/t8hVNy/RhXNChY7prOhUROnJSZ4AWO9xofQQZ36D/vgfORtNfIJ7Bp6WoYXS9rUkDdEa3/Hdk9
y+mNInZW/pDIP/vHaD4P28lgn8Z/4mCgPC5ZEkItKjc1u/pS+uTPLzUKjyKHPQkUmWbJuP3skbWu
F76Y5bKem9YkU469DojmeE/lIwpTNUjE5di5T1vzMK8y2sdkLLBpPeKoOkqvs/6r48TJuDXd3qrB
oauZpwmtAWSqvkh8An79d1KdSKbBsQuFoieN7GjJRYzosShL7/GzTZ+awAmdOrBvV3Q2L1bKoUj5
mWp3KAsjAOdJeH6n9CuQt8SE0WiIHgmVF+zCLZkOvgcPF1aRWAk6HCGaJupnjhKpBQlm5TCDoIOW
AStTJV5JQ1xSPCiKMUV9HrQeFqBg07ch/3WPANyVL1ThJGOkbFgml93AYLxEV8KbvVB9RCUqdDXD
zvVcHq4B//DV+SpmA5dQk/v7BLtFZO0HIHWhq8cT2RhByvJN8b823fkoB1W2/37ge7E3oc5I7i7T
62XRgo7rbGD2SrR/8jkCbzusolE+yxO/oEXkLx48hD9bzRnb39K8CPx3kUxQtys5jNR/VAGAbIcl
hU+JdE5cpKkpVFjQZVfOAwkOO3cnX3BPb3nf7I9lJy0p8u0h8W1dJvo6YlBxqlp1ZeKgxu+AhgE2
td1nI6ejOGPoystfsE4obKPaSlS/j6WMoi9GNmh0m+8gcFpRyUhSsSPJ5MEFsNsVRyxXDXRJ7qjk
bmAfqI38bKkkyyJvKTHB1aZSN45OJkWZNjFi4AI2a2fd5efPwNAorToqXLwRKYueU+wk07T/5J51
TBkrpXAqx20eXyPqm24grI9iexPN8bMbZrusA4zlS+IMIGjKStz1MHrtqsWfrmsNrjTu/LPsxlAk
ly9iXLtlMHYv6qVM8buBW65cvV6uGVMU9/Rdyd41BkM0C3u3DXF5PAh+JqmC+j+3db/4PW7fBIL9
ieVZ/k6CDCVwJUg+PjNNVyS7iwyyYRotKFCGxnwOae6+OkOagXXwpz/4HMI9wEYsKkBk0Gv5Il+H
3Nl0YM8IUZmArfCkOyoI4GDhBFTU0j22sc/2d99xLcYdAh1lMN7zqBbl90qmuNBRaLsfnf9XFr1h
pm6mb+VVtdpvRBWJ30bLnw1pVkMD6+Z4YK4uYtNtCtK+y8t17iZKmO+BYahHPLh61PTeRTZEHNGD
oes5FCnu02FXsRRevxnFnlcBkoWoGkrWKth/HvPWdLKtviXtBZEPaO/l3rgmE56MhB3ztsvsXFZ+
lUxxXBv6jGWKjP8MxjvclWXCcJ72Hk14CGaSz9bvagZtvGGWcmZSvCAmgmhMIWNOR4nKYp3mQnjS
AZYRoSbFg+9Z5scYNT1O2FPsHbmkEBdaTYSK0+3r+t6CYK3EPouvFH/hUsS6EnSdWV47vZJPBP9k
h/P/ppIh+IOrI/b5UkqjH+JGLWTU/Xak5I/3Oclzmn/YSjM8vx2N8Alv6x6/zJKyxPVf6h7PYRGZ
gkCTeTvF2A9gu2m6XUtdLZlHvIkVl0HLD2BSa0Qg6KesT1pXeaPFH04WE0AUNlzDUAx4Y8oRCoxn
LpscgltQbFvYPbrB9MTLzoS50r6JGtshcrBVpbLe8drbOgReS52WUxn5aCbumvQNc7Vqe3OMVEQM
EtAqLj76VhGFCJC3g6F+eGCBamUZAJ+5liFSeRZ1ciaZvj+QPoszNplY4iGysMXZttmze5no+d8F
LeQqsZOEDqo/gCqamwWs47xtpJZLoiYFKBHGK1ZCExV5+n5/eeAy46V8aRdGcHZXaLA4cyMRNonA
Kucnp7cxxB2eOuJf4I50K5+dyEPU48FYCdqtAA6fVbdzEcKJ7diG8yxbB5AjLMgQv/wpbQAAoG/u
un5hSElkSrE2O147VJukdRPuWEBs2TPJOk56yEltt2C5JdKN2REfuL1sZOr1dHSRLidSARR0303E
jodz53N/QQo6BbHIKpUzKZX1IunAV5WhDknl3Z3PAhRl1Mn6COfeaaUK2dS+4l6r52oQRziUMWG0
2i/xY8EVRIhE+nfSn/kYVxuV3gucHV+SoiSNqDMDeKc5PIOg9wtarpgj3fx6dynvaS9f4hh82rMp
Bvb77BfcqoTw/RAvGy8GWA68K1yaUPW12xE9aEokUfUEIFaQlAGOD8kr0kuQwiMSTNi98Bp6qO2B
hZbeqGcjgzlZ8SOqNdFRFLns62c0Skx/XLzhkUzlS3HkpSn/q2buhAdhU9omopR50fuCV6i5qI9r
wj7P5ulf++2ADVzU3GqpHjSFkMy97U/ej4RUormtKvqa/A8f6hTec+f0GLZOPiZlT1XLhkps8TER
tB3EHlmgJHHcxZ+hoEBFB5c6sExfFmvDHnvsi3ldTG+MTtRPXlMhqxcdj2QaQYwm+fTzJE711vzX
U2oXd1lrtlJdijSZzJcQv456OoOy5Hr6bZZQvZmQlDxvgADgN4JXiFv9Jum+4gAZwjHK317Zn3za
RK3CfZUOeuerlhcMb2A9tziAswDt7c9sj43wFQfBT+gD8gQE5PQGlctDQ8U2gU8PjbzxtXhda+Dq
yNOH5+d4shVNjHoAsA0CV+M462Ej7bcgzPG2s+07GVNDDBQNwi45pmDjQoV+MHp2dkg6gHMGFD83
nxseVZY2wYtD98aNdOqAQEH/lLB7M4DfoBEDkOfChGf+Sv2nG8npQNWrN7rD/f3XwSQIQYFiWaDn
76SuFYGVt9CQ7AQE+2KFwhlatlIwIONaZoPRqhBrG09LIhfX9z95SGXK94tJltgXnEyjtKdREknC
/qOkk7vzU9ExRAiI6RHOxTXa2qgAtKNSRCXqNePCytN97PIX62L0RNKKzjnLKGeKSOPzVgXRbGAY
V6rYYlQB9qqvKgh0Ncq9sHhJpVbzXBqvGku2+fo0DRE7ub5ZkawmXajEIpZ5fdkZtLNFHrX8M0MH
I18zpkiSyi/Ap0N2HEKa+hZRfO5GmdD566MTLs4x7mMRMObPoL9AohWo41wvyyQNvgk36Vq5weuA
rU2pGcGZZYkE1bAl2MxMES2kOji1DW4siTkDYXIntNWibnKLicvh/DK+tdnpDoPKVXlU7OA/w6JQ
nWmXH21fdvewzHjOqzl3W1vqjo/XtiGaLQe73m6Rn+pv4zxKRBs4eIp6mL8Sb9MhS/kX2M/4ifm1
pcZLvsCVJC3vYq3hwf/LOUeIG3fiD5aX5gVpI7hu+G5Br8WsM53txsh5Gp09fb9dKCVqeVDb3eja
3LO+mh/Wn6umyZuPdW0OACHoyaDrB3nKAGnd2xjBJZVzZdvsOtuQl37zYbXNF188K9yIRFVFwhPJ
hQ1tKYfD3nyJ8WkY4Pfz8XB+8/GRJc8E5l0cZ1gkXW8WpcnVLN8/CtmF3ReDYVVFdIzoaXpuPfxc
80QOuRVczWItS85V0jD7ZfQfaowKvNhiOm3lD+KgCzb8k91GQ/jYW0qvYMFaaai/X0TrSZDVJ8Oo
GwDKvDaFYDgMOGzyYTIxmYVZIOroEWC9Y8nf+JF9i2tCPZm+Hq+5uE2SxIs9/SsGEieANipVj0Bu
idQqm1KBIQ6bJvbxBfNHHs7VXTAFFxTFQpomxfPk+G9SEsAMFTKfGY8nncrbUnZfmMXDCoM2LVKc
D/iFXatneSxF89iBmqxQLDAky5t4U+AnKgm6w7LveylAXwyPZgNQeG8s4+Owi1IO+95RWHuqXKql
Kdz6sLWffl0FsXAAN75BSRPp+9FTTXeCqh6hY6ZtUWyswWeJ1jdOCK3B/yn6BqgQzp47WyRn6kK4
F62I9rS1YNrLBBtIwNwFHw08DQ88WkRFB6rptonhq75U5VrlCh9FUl9a5YA7Kslmb9stGcNnKr4c
KeiMZ2UzO56kA2zC3kW7dtBDzbWOJP1qngkyUrUDFFXgtvd8uXLgB1dqrHYBF1dgeksnjjmsQv7h
JL6oG3idjhaGmnQAS/OrmVvonFJSBtA7AMwUEw9IgtNVbyeoXwGSwqld9KIwmKLAx6oqEHLc8Htj
Emv2MAckHz73gUGnUZLc6PIYxUaJQ67V35SXzS2V+QF9bPJw7GldlwwazbK2iDzgU10IfDilds5l
CnYbYl1ykv9PzlHyRxDcup+vKMkLPhJV/HxDbmXA4pqKLpweJgPiaJ09mHIakJklm1W2P1heqmVZ
8MPs1cdsRWqzJR0P8ccbQ0+0L9Jd4CsU/rhu0zKtMyWC5XzsBNTPX6MzogFKfvHi5by77EMT+S3d
cUvWDU1rMQnXvzypVznWdhLbByZDr9pQrbqDlth/dMCDOAbaavDAUV7c30Nmm4D25LA8p3j2k0nA
tgSRiCZU1sDfsizi1injp1cpmAot2YuhS9gbk0RpW3fpylDnTde11Rr9pEvXbbVQ/ztB48TeVjB8
ZZBrmMdR8h/AmNtL2GAVikb/eS4C6pCfOqCoVolcy56lroqaN3yytiiLdAkwHpW1lMyfqgPy2wye
LWroZc/EchL9LPeSmVzlPxNfthYo+fjj7OiNWkRak9EMh+nXX/5L4WGsbh+Swssar4GpTwZhj1bO
c4ut5xh8wI/kQPHE65LKUiUBUXb/Mx03PRwr1zIfMj/2t4q0ZM9UOIzTvRDyeO8bYvt+rVusAal2
o234xf4Aaqd2bmI9S9nRSJ3Z5AGKC09KGDgXCFtChry3pHibYi5tJoA6E/owJpwqNVLBig/6ul4c
9ubY0lyI1p8WHmVjqijUYWWVQNBm6inbFqJYEU+sJ358/3xWnPrTc+5iQdHl6ma/8/7Ku63vYGwv
rejTMoKkgnjZ6V6lyd0uf6oX6iLu0d6g00OItF88FKFRWnhWNOrvCdJsHZWho0tU89w/H06Nmm+1
ZLgxwxKkGelCpCbvyNi7ECU4ZB9g2HkV+uiIWJVMVW0aeFboSHcwLGipAKxdolqrBqIPeKLMauQB
wfEWC+jn72AGw7StbGP6hZ44H9tWw7D7GhwLceUaxAc/A04ScyR6wMs/f74SECbjgzb1Z+Co2ta9
tVz3QtUsdMg4v6komy2Rlwq3bsV8IDW8klokhMgiW3DmrIFF4ePWmOF87R79boBvF3pq6VVKYPZo
eFYMV3WHztaRhe4zShRnU5YHQCRj6TUx0fpWtgfX1xOAfXKhOp7R6WhdbFvNMcv6EGr7/PVOJhbz
AkCkiaT2DnwxKwCT2rE/a1c0hrgsVH5LkLtwyxUcOU+HY5bIEmk7J49DMHdFlZpqEQ2GTyYjQ3yt
Lp5ZDSHB1rzhI87tLgzu4bHEktfMIRJlZ96DySXi6YdBDKTHhTOMyOvRO82F/V/qsFl0VXA+UvkX
lYSwJ3RDxxXslUSMqZhgs1zWGbgS/BzBJmy8kzptIgDMFeTBzlIqNkzYPDvAHR6D4M03PitsiCqx
Y9szWkyffItHDtc4gB7p9ZxlT58NlVF3nz1R1PCqY1doxHGCvnZkmLywjcgyP0/0cZZcR8up+GCB
xOb8CP6aNXhGLScVheA8PczsjFqPvfSCVKjpsgqWBQQJHpaoOHnvCusfiMCQNKeI6DV4P19vihYP
bsyuiUgI5injwSaubYXcXhUVNjxif78y39gjzLgCYbcbP2Z+cSpKSkML4b+julUMmFlbYoLLrDim
lxrOgNOuK6+N4aN4d9kjqwYs6VeZ2x65TuvQAYL/z1sSb6jcqVvgEajMo7rDd+vXa3vUEcsgLv84
+1Mp8M27oWVtPSPz9djWGTHuckRHBJRTqRWk9p6SO5TABWFOggDnYkLfMAXsULzadvFRaTN2Vu5p
kVxZ7oQ6fBDQk1X8LODxYHDax9a5XVtYovBpATHgpBxw9Ju3dwJthgOMCAxl/9CKLClMUOHqqPKt
sh2/020hIo/49aiwSe99MTQ/jgzFnyhiSwKlvXl1Hq0t62qAMDekjtWE1EO6PTriXzc7qtVADvON
Ti1j8veAfep3H2mwUVxq2g0DMvEGh+Qeu52CTn6wnjSExsV5r6flO0FXge3rFiYTuTiikUIVqGxx
FebutTigSpWP5BCb40tJmLoyNSYi8E72dOu7he9KM1jCXko8UnzLvYsoDN2hIxldsiYB95uOkeDA
E5imXyEWVm6haG3+1OvLNwm/MZwCXwcJHnZYxQdPKAYoaDSrWx27aUFJLW4WQwa8+/rbzNfLf/G+
mhrRH51oZ0sD8K7Fxuv7GYc1+tnoqd8+vQ9ycSd8l1KJUfq9ZhMb28krCTIPjrH2nDdrXhQYXTsC
piYMezpSLQlbS3RHGKdfNOlcz5DJ5HA0w547GRTwmfMh4zbZYChx+vhwnVk6l7p2J38+qYeG/yRx
cKPl6trl+4tMRRdbxDBy24e9vkeKHpEJ3NbB+Goa/34BZOWgfDeFHwVazy4mkaG7nzgChiii5jhR
KBluCTlhogjMU7A1Kl1SruKATXBhLBgMKxi2D8i4IR03P4+DxEYl/k710WoCJt50pX2fES9yCHhf
Vd9ghXDQl7DjvR++TMYHqgKH6gjDLCwsFec7gBspJ6HmdgyHBUnWbaYZylSvVRDzXvFybMs+1Cn9
qvnJIdGw0TXPA2NqhwwLPbOH2CNE/lSqbhbapCZOE8p2BHaWxr2BD7vT3Y1Ev3H8FLSg2akSNQW4
syN7ndCmVd7mitWpFRkKtd8DzizPaMyc0cjPbT2ncfiNCGL0SzKdxedXzU6XWV8I8Y+qUzw9qoF2
ziBubUZiS8ePsuwjcH9ZbwsT+WOUZyieDF2Tx30pYPeQDXOR2tM6rPu8I9lxalzLCMmy1N9ANljn
PbbjZFf25G1y6J2Z7jJ0h+o/FY0bc7dygiv3Lsa/D0/PHrRgkmC4HgP1VRoO22VYOLlqfsN2h0nl
n0Kyv7/DF14b+q5XbduQsEVEjJjAKbm3zcWSfw1gw0ZJRVykecVC6GWR2vS4ABvfYcGEAdpzxDve
HBpeHD3I8+MJh04TRyiQU2yvB85+XJ6mWcuR9i9T6yGwkerVGe3wpx5WDuki46Tb5v7uJmVUiQpC
VP9RRvDBYMkcENQ5TFAbo3C91JfKZ9tGNyFkabgokrx9hO2dGvDR90KyMLUAJ50myZe7TX/F4Unr
PcgJei29MPZACIcS8m4AzcOgcyTWiJtKc4LKLcK9U58N0wGCXhD9BvnMl0BGZlNiuYj6BoGKD1A/
0vkNK8/Nn7EcHlxidSMgvVVTeK4AdgdORUQbwECdHRKPf8BlCZ7qNX1um1qXJdODezT6O03chENi
H004uoPRu952qHeZaz7Vab56HYp9Ez2VUjNjoIVB0NbOSYe4OToFyutPASgUbYMxzf89difIcDM6
tVV9DW+x8VJn+PUQRHEZdHIYPgSQiWeFgcugo6oYdmwaOITQvtz2T0DE7urY1w/tnwP8td+//8NV
3cdsS+0A+CM0VDoPvuq55ZsWekI9P9TAs6q83EshN5oYNsApFazN+C4Qgvt4r4BMgOyyYAO8J/gc
Ij7N49YyCW+sFAaZWEcHHdrpcUMzYXO+/hHMNRQXSglERjX8IWA9Dx1ZluinWhaZujTCeCITJMqS
egTsYPvFh4EN5SbqDMzRNZQlDwIWC9j0s0c/wWJgYIfz/Sv34dVMXlSabnsslNsqN2fa2LO2rNDl
qjue9vFQqgD8mP6XHr0AHNMmXUBtY9d6zPCqIxnsBoPQn3UAwX1E0niBTz6IBVfHAylDssLsMEUY
QDKLeMnjt1wDKRT3ianFpOrEfsnIn04jqwvhYRsZ0ZC6Ew1WWWCiOrH9SgWPvP1wHXJOsRAB8HTW
sh2zAwt3W+SnlX9PufHJrlgwbOuq+IrQ9179N5KupBxAP8i2A9CiFX58N5M3jqmHt3qvWc9Y9KF3
Cp2JUI7CiH4RUht06d7jMwBjgPjr0rPYxRH3W33vc7TtDuy/BLjKpDr/RtRPY1aEMg65d81oqTo5
Wg5cFM+/8kV+NAxNf9gyvJDPrbw175a72+lrfIe2Vqcc9XfNF5MYh60itdclGbOJekFliqnWrT/x
+husJbbb9K/KlykXF4Z6sGz6PertAssfe7h7LnJZVOxAYPIqgYrLq2hCSmbnC2iNcBAhRCt3mS9d
zjZKtH3rZEfy09cZMjl/rXhbqj8I14TbK0rrV5u0ezUlc2wAsWdeCVuetbqdsQ8dr3CtSHLbjO/w
hf5XFVStJFDr5yxszM18yttG9TLOrAAehL7oUFviGsRuBnDp2HCM31ie76ogrom0LM6JBehKwyEV
Vmqd1eZ13BVrE1oBoSlqw6bhJyfCn63Cff9e/YVIkhWLhByTxeWV5xTgoPCLn+o+3f785xrPRnvo
G7jk50R+n5NBhN8NmazFm9WB29QBMaqq/buF03SnKi7JDn6Y4Ja0Nhe9PIBQiH88ep2JJkq3lJhB
Od5JY+eARPc5E/81BHxILlebQ+AaqqfpheQGTzFDVh4WFeaIZZ1R00PqDZY4zzliCxXselt4P1Ca
5379uytjaVR4B32LlE8VDOzxoOuuVr6/+4O9DkNKHJhgdwmXb54uSxE1d+HRuzRgBGAS5f/NVETY
l6ylMvfKahLehIQkAWmvzuhCXCcOWzFaqE2jwj4O/4x3iL94k6c/hlW6nKzJLQpPls0ye0Tc2AIP
TvVte/RmUsLBm+m/ock3BC84vgu/itfC5zY+kNXELyxE9MNqHlFBgdMDPJHOISOJciwqKi1xYQ1n
ww0nM4MKRaKOrX/9OvorYdnkSIWCmhABT5k4BHKmc+E2304yOFMIlp6edRDk6SOAf8mNjUkXPDFS
tRvNv48MGRdPPQec0VxRm56kY79vMnlCIC9B3nKVjGYVPO2Q+BG19FJdIfq6/TNvj80afdKq0zXY
4tlTdm8JgQ4Rugdeap3L+LzzYGd/5ae58cXZ9exAVYXVti2Mj33kZ8GN/ezyhIVUUadAB/HuPMDv
YFAUMZPnIvaAfKcix/TwVVQkprv4WYVzLIkCbvVY+nsT9eLNeVUlIQS/GTADf7iGNIi43nxgH/LD
jlZGf1adXAJAAChnHzkafA8HrpZaqSZr1gOuxwmpRgEUz3uAdeHms+j/uqnjY/pcr7zn+HQYfBmI
0McIeurSzk8ulhZcfl99A7qOu3E47pDUKuv3kyWrCsErZDmz27c/E546Gbbqv0PrrJpFpbooRghg
cfQ7nAokVi4mDrKPrAEq5/4iUL7HQOE+sStMJFUaeuqvlgPRdWBfqqMwZbkTpFtivFKuxPqB5QKU
I8BsM/ui7aXfMvC+SiWKCVkQkIfkUU2OYxZnlMAoPKw63wjcSLrDSAysrF4uIXLOU6zDNxesBPev
0dLAU/umVj/Bsa7It5LJnbQrKJV1SqYY73vIR0W0eFBW2CL2+KoTg0bjwe5TxZr0cnwZ1gEGkivP
cxPS+SNFDP/j/hzt6JZLEQAen4gTBYulITLDUVZ6fXzoYM1mpgWb7epvss1pGYg0AOMu42MIX04n
KfP6Jfr2JW0Z3VU9zdFwxyN/in4M/Q9OOwdvxhjsfo92c3oc7mUh/bjK1B3GoWGuRZ64dAT5OFny
LwxhDczyZOrYIrcCPqDy9LjYwOnOabwXvGO6S0gT8WS6ymBL+ExxMXFPqlNIH9hrQw4kVpDIpYPD
JpLB9mlgb01SzLJzHzNGDGtIYURxN7CZPlzDxMBnPNBtvrKwUvWIneR7ecmXkPxxKs6O6VS7S4EK
LzbNOdxfWxHSvXSNHLU1ZMttK9UBS3eXYRpyOvcv06HWDzPo0qGlYNThjO+BwJjYwZOzk9cecd37
ar7Jnj4MrG9dCD+xTpeokFP8U4yDaxG3C0gfGNRHQhuFJikqWPumNlg7NlLg93SGjoW7Db4imQDT
ZIi2RMyrtfDTZDrqhqTRVGeM9oEzLR1a6w/e6qAD1s0UItMlNGmEVEW3Pc3nycfjwFquxUs1hjne
ycxgBy5ZCjyyLupq4oiFXq6h/2J9q3WPt6Q0+WAECzbsfpp4LngBlyUs5zdAwbXcfNJP1O5UxNaT
8MLuMkB8bPtin0n/afGLZQfnJdr5dCcaMP77Kka+NQdteK6lMAQ22gl2DSuOxJtexjXiBJbejLiD
rDDzMp7PG4foXQV5em27Ud1yIL995TMOhgvyjStfv+/0dSIRB3iORltfcBsvarDegc1XX+AClHNy
AF19/C33Su+gwvJaF5NwNpcBMOwtm5YKOH0zMY795OrWCVp75zdnBBQ3slFuqt7FNGzVKsGe3+1H
ebB9YfwqpVKUm6rj9L+ddZk9y8pGb5A69HIiBqN1ypFXgTDbXrY0eG6nA5sCtj3te15fvhrqPEWZ
R+JV6cvltxzc2E8TiQ07U7iURk1lkIAI5AXDlH3ES29mdKixHROKq4+YH4bKjsgrGmjplkWvEhj4
ztVGHNBQXQS5O63Dj8wTuZhB4wbMFm8C5TL8BDUOjC2wWeT3AlogEgOunctLFFfAEzs9nKuqDyTe
0UeruuDli28o0Auj/LhSw3qcdIdHpifU4d9o7ztRp1v+2Ho77ou8Q9jbpnlFbwSMl1SMaT34Jxz5
34V0kCbdzXE+7Db66a94LtB8BofUtrOt5UdnyBsDYPWVxjtHh7T9QtdnhJ0G50pHWYouKDFs1WJq
JB8k1PImvurusYsSJQnvqRnTKHuiS5e+Kq7Zwaayelm0+7juzaDPZ6r4gi+iVO5T9qZTZcYBCNOf
z3xyYs5NOsx9fjsVY2ItdzC9cSWYdlMkW6h3ElyKzGuVJrFWhdNm/qi0LPOA9Rmo+ctMBUWYB8zf
fXbN6Oyy+uoPYnoiipbe1dmRw1zhn2lc3FU71jrLsj1V1Yvs0hypoSeBsaNvVQ++ERW4TqswB7lO
FhDgqmIzI7krhh4lqBOk+oZxNTMsZgLXPm2ujAKd5FlF75ubKH5T+B26oAETjRQ5nPZlZo/fiMlP
mFaj1lcMl5PVa3YSZTjzb8Plvep+2wX71E+4lO8j2hyqM35MG3iGIZA9WFtkVDrGFPYuo5wgJjGN
erBN6srZtXxoWvfi3MQZsPuBusTZ7s+fcGeb2gxNXDFuawL9nxDLumccpFiKayjpWS4i0GugFyHu
dcVKvaCk4SaXaVnIPU2TXV6XeuhJlQWIKu480HfLNFYjrVl4Ty4yM4+4PT9n5ItOHn3659mtcitD
X38F+zbq0kc+bj/2fJ5wv6Y0NmmS46C1Q1yJY1c5boX5iOA8o8Tl3n/TZ5vctGXJEIeVU+Ax7FOO
84ugd1ITCH3CF1nyY9YP5nAt53BiRG+lpHb0S/VAK5DMdiOYpZLtBsoKO+QMkdj21lHqdZCEw4pe
gjriWzpp7/VeiBfYNejQrv3OqLpQYF+vQGXNvAkyGQ7+ZDNedu6qcDQQSwR7Yk6dv4U19TR4V3Fr
4naxYY+AyVc2Drj3KWcDhFbWRwJxhT43FI0I/MaJ7sQV4xIFjWtMZqd6cfMx/6asbJWFJ9DEyaCs
sQO6xxTWP1RdxLAgGy4T6BQPdf1mmvV2+P2jrdDjvnmmpIQik8Msdy+PcpZJmbjcLSq0lM5/qPWe
p2g+twIYtkbgekyCKdUB6RZaqnH1ZcpbOplDHbG3ax4DpNnplyxNMB5wmdQH6G489b+AyKSkAKIP
g6xyNjWm3TuyOw1CPkpK9TISXpmJVTMVBiWF2Nn/KFeUyGJTYSALrXELCr6R4N6sPvZ7u2Z9ixMj
nZG6Y6wd2b1v5pqghCAFnz/DPTN1heFJ4VLG35r9VFmorDUAiMlPDx/Xec+0TQdU1BmwD7a/8f/h
X0AP7879SWYGelTxRLIQm8px4AolImY++2UMtqS7tgiMjObFAG+VJcYD/+pEu6eHlSjbdYa1mH+f
w+wPAO7QDfmkLo3+w3TA8eQf62ACoBE57zUe/b3yAeoaYvu4AW0xWkr7y6i0GAZbJ6r90LkM+EvV
BJ7o5N3NwXjPQV0RMBSqf0pDBfiY/UbpZX1tv1D9C3jz0sYjZOlAXbEhRrN3fB1/tOtLbWiiVffu
UHPd6rsN1znYzHeM+vUb0rbw9dv0FLmVn3+v85LxzTWy8YqcSexPH+Mf+c6glFt9W0x6JQD7qz0Z
seRnbnRj+WXICNgOJT1BOlzfvzLIni3CvV5bYvsSfHKcWw/o6HZhgQsEeMAHL7u77JYdYZuevICK
KDc7vkyzLhp54dpCiFGQ16PNsIaX4gJlbe1U1pDTCTpfD5pJhuT7tkXMYyTeKsVQ8hW8TgXA3Qbq
rGF4kg+q0ZB+1ZdbR7chY4ioa3CbQ/2H+9L/k7eMlvItya18medNbdcCGl/U6Izk47pBG59bLeEM
SB6N6d+JYrwQamVJdflmEdBIqrLuGlDh1QPRdlzKuCLEOgsv5rFSrtdAwwMuZTG5R/x66VsquLXY
9rB+TFYctOFatG+tRjkUMvewzG8rECEMLj5CQofP7aaRLImhCHob6DMOIZmZpUKScmCqZS6CcZdR
JgDVN8uTXedqjcVF1f59lhXVPwZChWb+klIL+5YL/SLUknF5YFSRjsX3oPSacJbb0l55o27lB+mu
dPtN8Wcaa8Ampe74+Tr58SbkwGZPhdBxdLET+Q0MX6G7B+fShvQqyq+puO8cOlewwCmqQg/ed94J
YwTlw7pDRlickhG6krdL1VoJuAvy3OpZWnmPEpK9OifHyB96Im4zCGsc+VQn3jhwDCNRFXglvK1c
hPslhEKMG2ytM+apsNt58k/BtnvWg7ErOd9aMZ4DnWUGnaFssdTa7U9cV1nTA++2EEQMt3pgNiFA
snfuZY1AzIyQGCkfQMcz/573eSjJ/nMn/oTG29BriMmgmKVx1ONQHGtiNe4bsU8nVR/WBXeeGZ2P
TgDxty3ydUIj7GU+lt2oI1p8797JFQWpnsZUTRMlWhN4W1PEdJF1f9RbeEjC3yTGZnMD9LSFRQEG
fjGai/rCojr8j1Bd5kiu2top+weevEwsvI9S18UigT/yEsOMNKsO4Q2dItBmVeh83jqvIsRrXPUI
gP3lYOwwyqUZ3Ge1/1P+haE4Rr/Sqp/kI1cwS48gPD3kz0JfNdwuxZZUTIDzJHj809HK6f31hP4e
i7LpjZ+L6srXtZ2ZlrCXLMN3k8uljThwGflZQDeRYEy58eHRYQxcccsDc1+gQoA7Ua5oWYgYPKIF
eL6sfvkHHAPIqRvWzC04WK0pgQTMNmc5TvUkmFOX3kHK2RcBkXtw96SCaJ4eamo1p/VIoPxJoUzG
py2yy1CNkM9H8hQdmZWyq2PhM+d0YQ9ZJBTHiTFaGYtUNnc7rKDpMKBvTSooigVWRUbTkkEwUCZs
LPKjZD9XZ6jb46mCPV+sz6/Yb/6FlooVzGSfiWY+xP2ks8W9sw4OIqq8k4VHsw4+U8wCJvJkm3sJ
WyvK6CjB7KjaWGg0vd4xFK+vfMSJOIEeehWag7fwdmkEAqc88Vexq8kikwHPBQnAZdgCXBcR2JhX
vBJqQsb5TvesIC/a7YkVqlBZBMU82CPvMoSL5crBdsdGkMLjmZwPbnL8nEg/s/cGn8cHF2SXq4e3
qk2URMFArsLvy2h6ti0CXEKlxDvmrsRDNULnMIqHwjz6XKAAyEf0s0LPomMw7ECyJ5gLF1Vl1BxD
aXNmnge+l41auGqKDSV4y2+vcoByI+Fq5m7FnA4vaNI2akIftKhNc2/9mpS5irKfQOpzdVXAS8tl
FxtokXiMNhZkMTil4Rl4M+v6LVZBCOpgleLoqh+blM9y/EEAisFn5knrljzzinhsjsYi2QT5N+Xr
Gy2vH5XXzNdc+DLVvRQhxu7r5aC1sQzD0IrLMDHufYHem3nrkpmtmZD01ugBXMrX/16s6QmgpvK9
aoWvjj/yp25tdzDxklZqW3Fr8NhmtI8D95cYt4gc3KCrrxv8uCThNAObDSOHe4gWGiVjrBsXvZMf
XPGssU/YYac+Pyt46Z348lq+X9w89Gx77uJQZDK3NuxVhza4ICW4/jjB5eLBT0IOzs33MoziMG52
UDTlUy77eGwyIDsCArwGuB22Cg/FzsOjDVeZoAENyYxZZ7L2Tj19XtBkkQKuEabI7HD8HPyRdftZ
cFBvixVObvpGZ4BgQWthqFdBO/ZyoCTHeYbmuA9jMCNNl2eQn1451qzmXrmwPZ4cQp6m5VgVOik2
JE4xEo+luHSXzSp+3gRjFmCsavxIc8xD3l2hf6tWbMqtLwosg6ihltB/Fw3T07zM3RhcducRYBtb
9ds28/ZrTDIusCXTMOO/OUpGvrtChqNqvz+GPe+/faMiuYmYUxoO3nRb0x848T0Jn6sQw1HV9i0w
Zu0qh9fA3mPtYq0uC2Zt5JF/6j6YhbSZGJX0oqICHH8GyQwXQPCmTXpVpmN+xmj9nupG5Vwahtag
z3N0KseSmi0K1keKQfBL9K+jFqGSXFVOOqd3bj9hGnZ6wIhy4mRGdJO+h5bjd8RttjesqX71Qwl/
DvqaVzp9ZqvXcpVXn3seZHII+fcxQYzdvXqfmWTFTk37aNc4xouBfderpjrftfcrM+1xNWetiYjX
v9TMW5iEQdjQRctMqh5Y4MwHRZD+KoYf5CphcPPUkgmSROzlYjvh2B4cPp7ns4Okld4mIRnQSbjx
NSJASkmTyrWhQ0b0q7aANOtYa1bOBd5VufEg1OeJ8uTSPMDPJmRtwkVggHbcJP7354LroQB5CsWt
LflCaaI+sSFQmHc1eOpuqLffDfbpdiAzCiLdcX79DufaqcJQWWlB2p8aDrZzC45q7JCIhaxSRLA5
RD8l99qWPmxxuKAa/8BVcERF5BLMhh/A70ERZn/fXsTTMQS0mXcPcIn6bVLTMyc/C+0DTyH53Bjg
Hy/mABV1ODWoajIUi3JJAPG5HcyB9Vka7Ek1Xwnu9Oyd5FSmTaVs/nT6dktXeQ3ucIHgrNMYidwV
od8t0RiS/67cu+gbHh0ukDPyMrU/hG3HEpIVAwFkJ9S3mxRkqgT+0YpWf3LZZWa8/hGDnleUdOS4
zvEeEUfNrHsHFLEhqFl54rYiaYt74ZmaUaNkZiXa1oGjhz1HRN5W/0zXRpuBKAfNI45woXf033QS
udiW3lExeVdcsBjGjRXJg927+Bix8cd02n6zZ80zviUH3l7PjyEbT9NKz1DcKmdFDsFwr5wO2MeL
0mNFqQJ+Waum1NsHF5YOrro/pFrvS+ONwhvRmZXC+w+1i0QymA2NZusvT5K9mCZj3WFzjlrgDlv3
5P5hdR6smTHfbisLVAY2RG4L0j/y+4mzue4VYQfXzvKlkditPu7wG/6IeeilcGuCS3bwchbUr8i8
UN6cQplG5bJGFi8fvJIZI1ljz55ZvXa1pBHL7eHU3VxBrjxINlAUN8aQkNstAhv91gjKnOZe1rjI
qrZg58RKnQceRby3y/iob1Q7/w5kCw0KgwMtxqI/idYVmcH88WjFdDlgBnXYrv4xWG05ZLc/bhh8
g4AHmxrRaM+YRtU1aDAM/YzBHuWYlkR4XiKs3UrRUBg2KEFKIRqLc8zWZe2g/urUEjHLz6GJEVcc
UPauJ8cH5DPl6HGnXAFOS7BB2P077I/PRv1RumABUr5Z6vkPMUtBRMM1G7G4igKJjWA0So2vSmJ9
60U/zTqW/0Filn6vitvyKzECaflGAUKfLVSz9r8YxipYdytBDHcBFfKQEWXO8niLUZkRovL2x7sC
diMrxgnYWKyY/eSJmi7O2ZUahPUeacYu5HkxLW6Eo80qMDke3CAObl2fW8DaX0UhIRv6BxYU2/We
aLY0QN4iUUGVRP533ehKNDB1OXfO/2zi1NWMaFkNnWwMaBXPbW5rnh09FmzmZCsV5WrwHzqDGvn9
Q77kNqWE59ifOhUW2Bjls/vfMetVGh1qzIxYM6PjJxn3OLhkC4vTgsf2of+6jGQxKH4bAlhEiJ1G
/wSqnQafP7U2q+oJ7MXc0vZd1c8O94lVz2L3XpS+qe0PezUJXo4tvOlVikWNPHq5PuLeGAbNWYrN
acl74z1CPKCUAEiIsXhPA+GjPd9k+K7eCnvcipR3I+nRa8s3vq4U0sEtBB/mFFltNfxcu4IQJ6CN
X/u7wQZJuk7k0i9pYVwGFuDcQDYdFGvroS3xsvY0d4MEE2RKs/QhyIbUaUizMsfgF+j3dE5HHXf/
IZzSiro8CL3bDRQeliEiUn7K36Q5rTsij5qvHhYYcJxiLY1TJ43IH2tBIUHGN1mzqIcv6uv/f6Fa
slXeuUK0PLoLnbTf7n9BpjsueOUT3DaJZLu1lLf16AmABGmvWKDx9uDqYVXMKv4eKFR6wafPa1WV
XxO1ANsczJIhfrY/1kPjN5IvVUsOkmfUoq7963Xxd2TQbjKNNbD7xSDr9wLvLP6gB7w1SUk6J/nM
tprEzrAB4Xpg7rJ97ynZ1GPb4NHfKqc79iylinZ/N1+macjJnmzuIN8BRm4jpp7aD7OksEPHpq7+
D39/dVZh4xR15qvhwV3mj2VnjYXn3gbyjTemTcZTXDLah0CPm3rbkycWxkuy7AcQHW28ErDtODdJ
QsVWqrMXi6XzhDcEEUGIlgS/uxI51NG4TCekeNeNGhnJ9sHKLrZnmbBvxz6F5SK4YNOyI+80nArV
UqvZT/k+8SzOdM9FNdNtGul+l/Mo+X43+pEPxYgj5BxK+/82FleiQ6dMx0UT01yIw461WfWgseK/
AlanjUtfZNRQmkHxWa7p9uCrLP67l2i/2mRNaNJEr4gmdfcApFGUU5iwvItJxEtKQOwHnsKLbRgy
vcMn3MtQEBQtXZ/z7MdEjSqfWuJPAmM8ukuhoFh7+RTZu0exYWOHFnGXM+7cuEZj/KgzJPRsygeA
OWQIqPxethPx61VP7L104ZJi4pkkTMoNGXvPkJ89ilXIpzyf9XYKh4zGjHqmoNdp1ols7bDXWuCb
IpJ83C3Wjm9t+qD4sM+NhYprm0N6a9NcTTymgIxaYGTvRbG2AfKlRFQvo3CXKkrYNPuCFZA3DbVp
Y0mUNLeHHwcOsWnJoNF4y34Q9gxdKKRlqSoPKUm2/mB9PszZA+kNimBfJlRDmXkQJe2Yk6sRJLBi
fcJokGL8cJGjiUTi8v9P2Vwam+4OzLXHublGSF3CRuUjDyl96u1NNXa0FBdpv21QXR50TfwgtJoF
ZKEIpiuVRg9+MdILE8ocgswVRRRF5p9OsSjoLQrWAk6BzTX9HajB6y4ySNk4x8aTs5V4Y3tXHlEL
ITXm/aWF59Mxl3KlZt9fJEMHg3dcRXZE9TKlQGGx1PAHPg2JfmcjOBHbDbN2XD1es7TVcEEJX3iy
JUFYGBNt0FQby5shBhFVA6guVhYwGk+0/aTQygm9ihPRhDVyY18HSs82tjiMpZM59eRSAW0BPkln
4CIjZ6n5mGZ+Na7brDGqLI7mokhE9EWHDjlBYEq5c+ulfwrWE08ecR9gE9gm5+Jz1VoBgZRroMZg
qKoBsQs03PoiyJO9pyj274C7dtQ6M0XbgNtlvZs7NiBoFPsvWgqMIdUuwshQ07Z7w7kInqd1Y6jX
/HdyC/0ry7yOsfNd/xoqrEkcgS8CMPCWHM8W54VIGjlVQ5fJ8La/OJy/7cHcXJa0MPO9XtRQ98mx
oEP9kAGKbG8iJfscOlXWVFClHONh9MZzvOlwkTVOKxqEHoCzTHtXO3fPQiK1VMW9FCerpa3c7Ofh
jKQQqRfk/J4U240xrxSE/5GkgGk54RVIRC7JbGDrAedOCJHzVaACIISTAXlevp21J5xynukdQ7j9
LfpFhy4LZfoPDwcPEu9l4v+cUBCPQyvoIY74mFOT9HWYkVskeFh/lZRmZJbtXAn/mhnBR6fZWNxA
pw19vXv4harcF6v1mgL6vm4HS/rJjTLQw8M17z2euf8Ls2mS7STgjDnk7tdrpunghyVjRLG3nrJA
kzmTM7tWPa95GKijhTyVMfeOOEyQumkFxS2CQoK3+dJazhZsSLl5zCEV/IaqpwDKTxPhggRyBJRz
+oZHh/jCqL6AoFJloTifH5F2P2yRBtVdTvVtvMqSM2BncaQLqPE6bCsWgpvHFpjCRlhSrvuCujFy
DOam6afh7xaKO+GBUbL3Akpr84c8W2W8noh/xMJnIBE+DXP01JD8pCj24DoCAst3CNLYBifivvmh
+cnIJP6vdEKULeY6JOt5BbeM+WLDiNfeo0xPDOs6xbt1XZJbiXSZUmZIiz+dwnE4L3UjAMwo+86c
pErt8kShrpzF1ajX9tWmq1sfMXv1mkRu2lzgpI3Inv2yDs6al4cIg3tJOzG0299SzT5XkMTBpZ1I
PncFXy9u0EKuwUDJkxbke5ew4cUmaNBDhuRCPbLDSxwMIo/6snt/gLqzRnpKk8OC/cx3XEHGONoc
e7bvgPeIBESexJD0yse3j1XE7NkMdhogLvca4VAjx22vI24lJvRLLZDpeCx1Uk/TawY39ejMydeK
5rM2wHX2HRC+yU0/y+N/fAcqvvgenuI+QTP6yl4fS3s2U2DhltFsXPU9wRxA/XTNGIl0Sg8Mukxf
s9qSppkG0zQ+OyXIxzhF6GTioVmiFc9s7qq8VQOovNn5W+xGY5LAyk+Mtum0pw3wSACW4up40YbW
CcDHBX9k4fwNvDaAT72RZfHXVj31xpmD+JY9WVLnwqjhK60M9tjIY2chq3h0pJVqQfsZ9MTibIas
G4nePzxJTQGCJtcd0vfJgbA0jYg7tOoaRJXNTbIJkfTB1dMNKj3dnWlMn8bVVrQUygMcMtlui5R7
whpL8MoKBPBbqgyNT9eAi0kad54/Lkw+dNUjK05pHjR2neh+UlWTOWmlFPIANUOaZSUZNp8KIcOX
Ptns17L2hdTuDz4o2X7BhblvOhcE0CKUUMoJHExkLlqjEcbg9tM0A2RUO/yqNjFBRXIByA+FlNX0
Ds5rW69u/WNg0j1yHMP4WHkmug3iP+fOk5sP2NvmHIPjeTfcKL+RlaFg9EGdia2Vdagj+XzwUiOb
JkUvaWPiCKM41R/qm/GnSI6qI8NwoHmGd3s2qPPAWVGds/KCWV26TGUKWcibYjQIz5ueOOZb0fKR
1MQElhnoI9ZLwREmjNQRHg32qWNZFRlgjwuPBUD8BYZmxmPIO3cwGXLghuXoZwrPRFpLpEv1ZRql
4Jtr3bT71UA8TrCEiZXUrVjAc855CqQbbe1iAwSSsuDxWvftzo0+wvvHDUsXqPfHD1nNsygHyqrn
4RzVHNV6/dHljkK7wD8Fj5U6+5tjXlB37KJVKz5TpNnBlWX0MikNwqatnfXlg9TNi4BtHp+FS276
YnAIA2Evadu1uFlpZGMltxAedGMtH8VT3DE0EGIHPG4cpOyru88DEl4YvNXkr00a5QgJTsztFohu
oI57tFLIf+eF3Ecf1VEHDV+z/Fegoo22P5IuoX/m1+5hzCqDoBYSO6rbRBqg0GKflDBLtScqx17b
jAFOf2O4QnKyEQmIFnDGurx+BhR8qzh53si/K8OzRcdhPqHnUxGOMxuZETyeR0ASH23/Nsw6T/R2
jVqZzVn2ytEU+GALXqDPdOMo4IMuxvXny6KOBbZOAl2eBlYPoXjg91rdqszEqT7FUOHwe6NIyct+
PEoPX9vtS+In5mOaNl/iRRYksnuc2fKbp+BQC8Tl7ZFXdiB+xT7K6K164SKIWOYK/hRJ1f8Yn3Cq
6JKG6DVIbU1RhjL9M+cU/9AmGIy5cfsD1X7x2Q2LTNy8ODXD4JEZsY981XZJ3Rj8LaD0SXs9RMtz
yZ5Okkd5V6UvptEsyfjUjwsCqjb/H1vpKG4nhO6Gl7O8AU2V4s4h2oV5FjvL0eGfCn8dE1rJFpXy
Sw6lCfPnjozBlY+Qz8HKr8DLJuHZx3OPdB3WXDU6YoGCx4tX9ipMxwe1xhWaUe12sr36O7sv2Gsr
Ko6fcrer3wM3T9bgHN22j04WoHxv7FME8/jIPNBJeWkuSZEvC3HpqfbGp18MdrjVnTC8+CGk/IKp
GN58XJ9RFoeu7tCB3OnbuAVI2eyYyg/1jn5ZE+qmoyE8ckT23i8bgrDlW8VbP+/aaFVcHXmFnTke
hpWeGGYglgFujz8t/AqUCAf7th1zpEk2Tx26tafPq0bxPhn9rxVjoZVfV8DYp6KFVxaU0823QGHr
XHSJHwxFCXx5ChGt5NcJ0FFbQRF+cIRHw8Zm8uCeTuiPqTP1cinhS3/LQ0LfpuuT2pgXHoUR42fI
wPpeVo9pvtk07fFMSyho8UKKaOEWZ97F5BuTlSgktTuZyp9IFK5gHHzOTgLj5LIt50Uzfu7UVn2H
HQ5MzgSXIkUVtJ19bl+8WMdXiZR3ycev2WTHAYdLyF8jPIG6RMytoBnCdRE1kLJYnCXKQT6Witt+
OgnC5UvWLZV+clWK0b90sWGeDEFPDpNqu4unuEn2axPLCbgj+K9uDMh7NFNn4rqZbk6zrJKiWRLv
mAojvDA1JaU/zVWoooFiXUlN3utqZjWjrAf1i/FsO5upsz7FWm6BAq5ciFzAv9BZriuJPzFcY+/P
XE9WoQ0PwkkYkFBOwn15v/yGBRlxxJqrQjd5yqmq73UOQbkP4KLpHR2vNxKKEPZz3nDUxPV0Uurp
rgaQOmDU+5/RCzKwKZ0WBpStqxGETYFo9/hnIYMcErEMjJhkxjV6cJcLXnxsZ72i/QiQvwTM7Grb
4H0oJSdyzrXVwOom8WLucKWfez9l1hnH7xtKBark0Jyfkz+mQaA//Rc640k8QwxXjeqqWhmjBMSn
502uswOl17bD3SI70k44SGxsG/q7zX6EwUed8TdE5myogssopkgzgVxQIdOLrgoK9RFe3p/N/ZqJ
RcTp+xe290Ak7VAFVr4ygLSeVHpjUUR46B6QuukRci2cw6aQCWeZ5CBfoS5Siz92fIxWjLNfzSUY
wvHzViNkuwNW8FClLXQ5F4OJhEdeW0YarcCB3H7BE14BR7nBu3/ExbLjn96PZfi1EupLi8ozhp1f
fgHaT9ZzZ5aXs/bc8GEILIpHizRhYrydHpS0csAXMHV79Ff9FNwi8f1A4x3b0N6xOsdpwyE22P4P
iwnEoxttae5oNcj8Smz9g0Gxa0iGSyHEudxeBnmKxapCj4YMuG5AqNs/Eosy5icZ0VocF68Tv4JR
fRSq0cho6RYrROIzw5G7P4C5e1Y+lMt1RMkoKcyzzka1wdKyMvABERmL7wQbzoTbzu5qqnipUcyR
dDjIIA0N0mPdtF4PlcH7ov/FE+Mf5tWrBHlilsWONM6mPl14n6nc/Zwf3cawxSv0m6mFg88kie9A
cBlNxqA8x5iaGY6xPVFywjxkZxhA2TK56ysxg+LeACjNnCKBy+DTz1lFlOvolp7SG2a3H86uMZ7G
UVf+k/kPSPk0MJCDoURjMjl5G9OIDMATupWo8c1nXncTAkD/0BLCXolcRvjgzraZK33hfDxf2vxB
Fxx3mtvqsqHJXuf1PAU0Oky3eOJi33i/NijUbG/6iQmCsbBfS1FIx5CbRlUsyqFQVDNZLJt1AWg7
8YDGdAxo1Hltd87ev3be4YqqcFibUYfSbHNPUmei7gVTGUuUDktxDW8mbCLWt1Y/sTw6lHHWTYgJ
9ZNZtMGxFzwYS/yg6SBGtE7giMc3UKy8BOXPbEC8ow66e2tSfB5ksPIqHeRsCrQ0Eb5Jm5OL6+de
j0RE/1BrJ7UjahDWfSBL4O7T9tkEOU2ViRig+ERZbdjWoV0dINXa5+YJWLrZDwKVeaiHLPmOPHJR
IvhZndFTY0w3JCvZgHWtrAYmLtqWyegSnT19hjbJD/NbWavG13Ogrs8UfrORFcwxl49U+Y389odh
OehZtDwqzkL1kUU3jJJmJOTOPCffktugyPmwPC/J49BrQa0uBFhoMJjJPEjxCbxZGOF1lalFE0RY
HqdxWGePDXhY4ywXjfCN9B37cQ6lpgX4lis5PNk4UHWjlw624HxPFl3+mrO/W//f5lX/6xqvZjLG
bL1JVGLZRaYdilVyk3ShIaU591L/PlWM8nGmX1sWyTqHG4rc4gnYkftiEqD76SzJhv7X5PgI1Fj2
oxS/LRhxf15MOKjGbVGNSiXoWaAH9n/pRSyYEhP7pBUx5ZKMpTDkhXJq2DAG9bdZvQDhjGDY0I9f
JxskVF8UP/4DzMBZL3OTiIvbTqFsVsSJkl5Pdfb+7oCZEubbzbJR70b4sZ0kSs3VbQdJ5Y/91pYQ
P7MpICLeqLi//1zBmrGDKMDP3hWogtAMdgFmzCYTTt1VMx/TeEv0nP5ZW9+f55S6X+1sBEAibWUQ
Xy1+rYytuqDpG3katZXSGEl5NweQYboafA7rKf6zT+sqw16ukbB0Sf/LO+C6/rYv73DIvpKa8o2K
kih0NBdZDCbH8sz0WHu2F3jTXWaOKk+L3ODBbBOrUq6HEwwJM9KR7RvjamyoaFdoRrIinzRtXfat
DRfb4KeI3qErIvNeK4aaetRmc2rRATp8o4mH9ELjnGH6Y917bbSIlhyGZF+3lf7Pc0KcggZN5wug
I9l6H//hfAw4z1tCX2SX0eAQrhaLdUww18SF+db1vCeu4Z5+8frlmNfl2yFx0JFIAT75yrQ3/RPV
6Idcp1ufO2MGsScbCpDeA+Gk4z6MZQFlnzx4RvuhDw4uHGb1LAWgl043dK8SmeYLNuGR8EBl9nyz
5qaiRzBHtRIkPyL0wfS+DBPoSjdkF4GxlEi/bCojO/lBe0i0jNIFZMDQcDb08ztIyxNv4yJmE5vX
rnfQuVrvz7IHSWdMB16PqhfWPHhOaIQn6LRnbQ4bP7VOe6wHGQa29OQ3axn9nHL1K3dG2BytDKMH
1zDzq7mRNBfuAn2djtCSuQQ6u/VhWoISEH+4YHW2lnAipi0BIQ/Jx/k9TopDPFXSnOkMcCX39tm1
pbLkWLX5/FsGokO8uMe+1AuwjBJ0nRJ3DJPNIacMEgVeOrs32qPg4HC9Q05sUGryg2ngR3G8Yukm
ENomF0xj+RvmXe49KpKvnEGs7L64IAZABFNxOgwSWdp2tIqy6k3rxnWX0Cwy0sC7v8Tt7f8aOYAJ
K0ZrBddf0RYDyoUz/aFXdOfgxIoZxuS0+cNuqChjTZix4jC0Yc6/XPN/zwv1jJdkiutXc9pHvuA9
DXe93vLA3nFvQjg16A58MG5BVyzhZyl8TTwYj3ACvFPgwyjP9ZyZRx5mxDycfMU7UNK4iNpj5pwI
Fl+EqL3+hWxzTTbs2OGlA4J2LFjv1rHpG+zzBsDLlDamzoNnuzG/5gLs8QW0/ui7PPxDtUEXvhKO
hBUv8bkqRY4gVXVfaBN7JONc7IBBF26AgJuFFFKrnyIpCWhGX8mLKrdOXpU75gdoiSJqMdzyp7ZM
YACDDLoqeY/bL3/fScwWWOQpmyx7E+KVWEFAIYvIqMkOyJ43tUrMdL3vDKCRvUZ0PytpPJ/+mwLO
AoJD1ssKNECFwDPnMPO/P8jDd7XYZjXzQV3+r6nKXewzpqP0EbK6tF8UW5j4TzTr6qN31BNPiWBx
NRPGryjV6zPGgHkh/thCQm62+X/9s2c0XaJP6gtseGP7H6ErVDLimrPcPkL/VwmhQ6P3HVOLDYgB
K29+9RY5KIMYdwuW+24JTjG1jD7cXf6R91f3naA/cW/QNeQ1VIv8p5hGaJ8CAqF7HioF71Fe4q6n
qZStV8zjQf/MYoEWLCDMKXcRxKsBAGM0va06/YRE8j+UgK+V+QOCVw5HT1mXr3sJK377ZzAqMeLS
M7AelsS+zpgTtYbt5hmrO+cWkmPbFSyYvByMYFuu8fyAeRTayGjX0CJgTOooU3BO15OJfciEfZBc
sqRFyqqqghmR4MqlFJpSSv2+cUkoC+bNS/pBBKCt+NYNUO9mReb/U/vIkbUR1lg3lmpoQt1zt5Po
H+Z9tnW2F/ab7FXVfx1KSM8dGjkErWaSpIQ5KyKhCChoFnpM0r+5qUiqQ+Kxz8d2xHV8tgMYpkHb
znv9eyIaQyVb6UhqUHFuY3gLcryKkk8olHbJ1KWx50vTV/Js0i0LVOZuVLViB0R/TXQfd2n73IkN
AbKGaecDIHWPxTdKL0c/fj4aKqK1RiZDv3l4KrsrMIfG4YINO3xSpoUB/QVTTp/6GcWub03yXnKJ
uWO3LDTXQycI2eUQcv+/ts63cUpnCJ6CZIZWUBqIlo7QfM3MUt10e3vRpjLycVdUnnr+l5wj/yeq
R9qDdk+1CxXhTmktidyrvnj6mSByX/2ky+UFbWYHsnv1wgbLP9Zl/z7jj1/95cFIAtapBfIm1QPb
qCUd66e2g4d0Q7Dyr/5iSSUvWdVXebE3FhsrEaffdcYmdUzmu4PAKbokUycJiR53mcnpVAmFex9M
VYz3LLXmhimpYy+rmFaGfpNt5fzzdHi0ket8taLwP5XM4G93QNuZuCUcXQI3OY7O9vBBtWurfH4O
EWUunEMedl8GmDH//YSMrxHHuCTTx6zSIv0q9fs1d4HrORoLfdnYtpmJz5oSwBOBY3V+StsE8gHo
DPcF21aGw3pylU455Z4YS6VLQIrpRcdr251QABtmnz9sZg73LOWhGeyv21+GmGl8aiCzOmcrraIG
7edHFX3leWlUe+MRc5SLVZaRk0kauQnJrQzyXasVncX1Ih+7m5GornM4c1EtkjN/bq/Qj92kXfw+
I+lGv8OUDO66yr9NyMxRXjex6234sWdrtoH3eWMiJ/O3k8iRyaLwB4EL3GcbYoHlyLS9XJ72+7g9
FN7JXK60oJmaSfXpk+jZKZG1i+uHuTdHhFbzVUgpUYuXN6B9qRmvc6F/s1wm3jO8FVjfy3xBJ5cI
HxQrw8X4Aq/QHF4m21FRi1vYwXygITcBPbCR5blTMEJykLqzayB5yswY55l5HMOsyt3sNAXKbUJC
SjSu8M/ZhGyfA8L6JIn9ga0wJb2FKrWwDJslWqUiIUf/rIi9wtu8v//CIEb84QedPPPzQILnQs9K
cZOhIE+ibZUeVnQUESF2bdGxnUBTWerHb2nwYyYwMFOoSL9ylMifxQRnnzEi22FRfpdjXI35W3sb
w/6L21Z9e5hj5fDCKz6RAvMN6NwAB6OiBPPF8xZMLcTdD7f7Sg2d+sLMblQqdP/KCDKFdwjsVpqX
rTWXavVPxnfTbsYuPm7U+0Mj8z0qtGrbR1W3TqBK07ZnRhHTjdcte+BV09ZEcUpkE5awr/bOQmW5
+E5Mllj0c90fxOU47iZc7fZGcbUggNDEwYonP9I6Bz38Khk5N8GRvf8CaPpVECpvSmN0MShQlJ4i
4ZiNftu43xHI3CPbFUeo+on1XbRmTd2Nt+dmTUXGRLfVw8S6Fk4Tx0U3oBYVs9grp8PuPrzp0lMv
E+jRyJ3kDeiQHhzOnwz8E+zcsXYZM2HERupcrnMHYBWoQDnKrz5thGsg59BmSJBZtrQX3laSqKXP
ofW+T/6L6Ob8J4dTivRnLAiF26F/TqCM0eWAVbKU5dYNhWIBL4VuITtUrVMLpT8jta5ELecHFsrA
t/0EYaG3Ysm2bE3vv9UeQgGGkHMP9mN4BASRazXlljBsJ8kNdDSHER9JXiVlELvw2ULBZZN9xMEd
AXHGUsVITT7nFxAv1UlgFzKPr6AuzAgOOwn7iT0j5NFHTMfSp+QTzD0jS6R7p6RKeceKgvOdedbe
MR1SKqJjA0PR3rd0O57D002DSZmP0PAP6sGCHctbpYzGp7WkfLbnQeIOmll7I7fxjtBVHNpJVw7P
WQ1p6h7Oo4VXFiQVMSNzVb8NTtnfvL4h3Jv88tuuf5IaKb802D9QSDPWfhwxoU8hmMjqco4KYL1K
ECBJWYQdGQ8Zv7yX7oZjrutfBj0T6PzJ4bRXT1bSFaMXBgpuiIuLCtvzBVkDWkxtUEfKklz9J2w7
kook4+tTMVgMwCYkkXqQZOqjh2W0j92bDZNMipdU1KX0u5iC2sk4Ro6CBD56mM26aaIFMR6PLsPJ
2D0fLgaegg1P47JkZ9jgownFO0LxZfCbmvkIlulsrE7YzjViyLRn0KwN44M77kOvOTphEwhS+j0j
61QA7AoudoWbjyZFETbjCIuHnmzyNIYkxeln4pSvFSZJ5prjG5LGXjPlaqQxaibvDuzxhmwW1IEP
3eEq//VZ0iZJZkZctiRjnj+r4LByZkdkaTnpAYf1pn6hSe4emEJ6haJXMAr2aAcIUuMCZ+hFwOha
ukEl4/xaV+Fb419nsnK2BqpBxwu9pCrf/+CNi6VKlm+CqedlejTaJuzkrB27lNhmF0/5TDQlQWxE
pOTuXJyAVi0b3aUf9JOFBR7+IxC19xKhYqDZH2IlQnLANwzBv6oy4YBVX4jnvUnt94gkgQTgbZFv
VGPRDsV+h6tquND7SPr8S8Lf5kEw6t+iCZkvlO/ipRg348gRUsXF02QFGfeLul3yGWmeITHjYpPF
3OoVTOVjXpvNrtUGPRM+ebowrW8X9FHeAUGRpm7UmNk7jAMnnZL+sCmV2DkhzXu5AQWqj1kWHtks
0cjtjKbC5kF2GZexw9D9G3rYShUowsISZi/SzKcAhKNaipnYqOXLvjpGuis0SDaq5NIcALthG3wU
XBXZRitydBxBeD5zOq+NN9gqCELEPqIaoJiTs70uZimSLS2cySgtCiaR/DMSLElbdskJ6gw/Jzny
fii5wolf6WLLwWkwoalZLtoZnvjQnw0EH5c5+WeK5eYe3rA2lSm2Gu+82Zke/DHH9aJYewuZeilg
s4kQqLyqFvZ9SfNDEueKcHeaY7eWDN4frXuEjrGlP/pzXrO5Cub6/wAUsTORPNTsRFzWSDJioqpm
ZaOaN30fjMtUIGbyAYqIjp2wob5eDXxiAz0RQcmNMN8VdESl09R66afv5nhoOQdckAFrZLwMYjQv
sjCTKd8nO/9yhJo8DwO5wSiPT0QYmt+C1fMSG5muLhD4t/5V9+OFu+fZ2mKEVgpiOuLHxQf00iWv
ab5ukPb06jzwVV2FvyJZryGjL7P1xzU8DP5v8gR0u0/8dykrVvxm2ztcigjVJyQFt4JcFZ9dq4YG
khC7rczZ0lAGUq8zRSdLsGo6Hnh9twPwYWKB8MfwrQmAv4Xf/VISNuBt73LvudvUUCWSoNlAMjnS
udm4lQilhdy7KMqBzTeWgKIKSR8PNwLIC58layUO2FX/A4amCmItVDQtP+FZ1FMaewX5f9ebtOsz
n3ufrYGWHd9R8EI3QK9iB5/8XHi+tnMt0dnu6cLKLfe9LFZceNh5hiApkQ7IMkXECgoMexOTMdTC
QusKblpuNqpBcvHqK9R7y+2HUDp9Fe6+pE8JjTV1JnPjGpeWordI/m8dRRRBv4I7R0fKFJTSZmWk
y4V+/dPLhIGWJ9kxo6JN5qny1BWCxZ+mJHXcFFKChRLMOmDCJ19UDSVCoYlz52ECC8FYXqFGLkBS
OltIYzSZlVePUuZKxLZgULQdL6yBcJpdPSJmxEvOOLmOdIWnvF38YSnYDf14zMtFw3xPLu4Uu6O6
cA8NHu7mYIBGwzxwHleh3TTsJ64qnn2JY3nBUHmpTJ+JtiQLcFaee704j7ISpypQBacHC4bOCtbm
wHnttyqBWUc7qcHEzIsrUk25VMNL+g1njg4TGn5ZtEWxY6mMOElw4Gz0f9LseWzAlWwC32yQC7FC
4DdHxGMCIlk0NcnvnKZvM5DvrP8cvDHNzD+GmNz2YyPmnZ/dklOFrtdbgNj5yH2+7onV4nTdDAcz
kkrJZFt8UM9ezFGZBCKXRT8NwuwMD/co8cuW8FmMrgie5hRg6iAI81sa56DfedrPSEc+sL2cUQkc
JYyAV/s5T+5mAdN4y1SkK3JmYZOO69e0LD/7SsxP/k5iLAL7ML1OUQASQHhUPdUPfLi6KGMDVTGm
xFb6yGru3knVlTaJrVqsOoeEb5g7eH9p6ocoghs9HCBcIksQ+Mu/9FuuSzr4LP13JuVBXA8Dp5rC
HiMDwMEgyqcfKBtyRvo5Jtnk24GYIMkAmQirV6+R8Fc4VWDruMWawFGnz91x68wDj5sjxR/3OCdd
GWzznOph8fyk4r07ze2EVn4fDwjNgLwpOPBsjh8Kwt3Vvhu0ut2qsf8t4na7/gCLF1nKjFiRXb+C
BTaZXJLnheY/dLby4Hx7U/p3MFDKYpeaIveYP+k0nRt3jQ0qjVnloY+OeLR73US99ivpe9L9eP5q
T0KYt/YWfwaSVQHvM8G1u5iPcHOgAEXzKe+vXYxHZVyXIpiXeRPTvbPgWWhxWhBz+xCA3llIrU30
1OXYFSCHXCCroAkwGaJAKKox0ye/1XoJuuMf7V6f2gRSRUQ5egtuBZ5+z09GtK2rx/jUjZKR4BqR
WWicujGMBg0yBpzBA0XsYUThDy15Vv9//IUaz1m1kCKfkP079tjLdRXbO2MFlZu0V4K4eB1WaSEf
O4JJ7PJXrpAP9Z6A0oh2vlBGKUtb5z8DFhFidvGQrvQZwl6rAscM5Km73KkivL6vn23IJVpWU8V2
ZbYIjrkhq1Cs80H1f/fE9WncC40VlKLWB8hwNK610sS1ZLFxMxFIQqv34lOBBfwpfn2oNNEDC+qo
vjddxjA9FZ+1dt1yQJrTlJNZFh5v3qifo9+B3xtzAxKxolryRFrHk0WTUDb7Q/LZk9i57aK4+N+Q
9oUM+2iQx5SdMUkCRY3ErsYQ2eot6Sq2bL0xo/AfJDBEz/YaSd3FkJa4paleTLGpmOJbl/x843sM
fNGLm9WW1ijrGXRxIJaC1lQi796wYymVWD7Uz1uIT7onM00LRy7tft06gHZMl37dfGrBPbedf0V9
0ztsD3BwlEnpyT578GbysZNlvRQjUH8MJNEzNNkSstuM5r0nKbynJ3tGW/hwwD7Id8udaG99ksNi
EVMsbIP/hDndac6Yyt+L9Wt6savpnGxqs4GpNVu2VN+k71hJPTQ0vgSYL3zIEOT91LRv9YIA2WiU
87hseCIt0/4VaYyfccD8Jq0JkFENdZyjSfiRaRnmj3gqJJeq43SqvY7nLMAJwuF94lwAm/WEcVTk
c053TBnONAesmwZ0TvN1G33RFKiAChAl2SVdV0c0oRe67nbfpDKJf1+KFMKhj6qoZaKHZsRou96p
jNEDi0qIuYZHVlsPLCZG+FrN6qUNBToTiBWFdyRV+YbOZ8yJSXKzwOALh0orc2K5RJVxQA4OfHjT
idEiJnAPEPN/6KqfBr6tLqTXZGjgyJZopVn2n4/S38ZaPDpHijBMu3xkm2T/tBjhgMeWSnpmoRm5
wpuTTA2SKrp3m1oiMeg92z6VfEcLQ9HVG8I3dtbyWVxog1vuCvE/RBDJZNiCssUTcaRIER4v8BBj
Ll+732SyXoF0zarvbKZBn64ij1glkdoW+mxKL/XT4Bs2klZ3NVlNBYE9qPj3fmRVwcB9UL0ZLwGS
BDONkIjps5SjQNx4PMkdBdOwRvSG00tI9nMbnld4v1MxpbqSAQqu5bfGUNX7gp5QoTVWu78HXzGq
phiGn9VLGfTzM8qqoUkDqq9lGWl9cQPmCmnsw6UlfpvKxzQIsrZK83ia4Qp80f4Sj4QOTpZARouV
Cc1TWgUEf8DjcfOa3X0Q0efh0RWQ32oCOQ3qzYvtlmy+3YBJv4ZMO7Y8oc5vpzvu4xiRx5qvBDsg
aWwsqPqWNCp+O69fCMUYCY12SGGvEW6Z4AARA1txCw5FxWhB1edWRX5uVM/uKGqrZKcl5z0wpE0n
iDs6s6Fp7uCV3VhqWt66O9D2v4ZV+6s2aTOMeNyFZ/s8LyYrICbtmjXLEtddHakD5L162+TNQuAE
jaDmnqjjvcPTXenI18KhreiyX5q0H22lapksMN0w/nY/DRWXrKuYG64bVjocIOmQK/xfVzGK0HoP
sdwHtbApI6Ex104evvlJec7fkTmvzVecZPhOfJw23Gbh14lgBadnZ4FXY/EaST4v4KE2uWu8G/wy
q7bzU1v4l/z9of9mtHcsl5R1rNNFDpgb6qTbTiD5D7fR997nkTcABu6o2TMAdMjSqAvdxGSNwYTt
ZPyUtbfqnZmbyDMUwaKqdFG3f+wnMDfP2oHrd8jvcVuWMULlD9VdoL1hFf0jWbyO8wxy7u9QaO9T
DNj8L4zSIGFpbSdptJWclbsJA26nywxKB9Kvj5deYyxO/ahCxGFehU8Iak+fXc/K/42RtFMeFGBc
fetAXrOWeeuPat4MaJuHVLNJjweeMJtEXZC8HE7hCo74q8mwYT+MIy1juSYmTUFjZTwZPTfDq1z/
6p3J4qcEnoh5jtbHWrpKksSnsseylNpXDgF/8oEJZm+2lPCFE6mevdS7uPiIuO7sGF12CVd5AsaB
RbuyGlBxpgfupGTYwVZiosLmOQECnBeieD0ltO8kEIZMirU0J3/oT+9L1AND+u2E80/5kPUFxTI9
y64HqOsodwI89O8OJD6xFIXojK7bvQbXvmPPuVRpl1R12Yh69YMPZBqornrM2Fq8YlQuzTaWS5wl
viI+F/7/ThCGbWaHbv1HCi2rp0hZwPqvtPgk6Hf8Pthj2xUY3vqtkr2cieuQ3VZTzp6d6lvPEAO2
r1AdLHrpJ7fOyO4Ej+kKI0gy4QQJaBVqAN3FwyLQB7QgyuY4esZGV4Lfr/F/4KBKEU1VDQtThI1W
oQ/NkBIbALfiejkWtLXHPVHovMuLeGToKhWEfWYAchsFFka2Jam41h2qifvQYRilmD+oQFVKbBWA
3rm58dfou78NELtg38fS24DxEpTFkIqpeC2vddnkP5diW3MzFF7C+/hVnVMM28FM+DTlrgpilBfJ
96k3FxZPp8WCbtkf2VbjRnp7CBSxQn1q1Bl01/fQH+NPAu/L5pqXniNsFpPI3w24Ux6Jgg9vmIoC
/JveotoyqR9fhJVEN3/vBPI4QU9F46NOb3RxLa5i+VOAaltBOTU+FE5NgcjtYOsPxtCcvdmFf2rS
8cEZNzJIbhiMMRj1PJ5/6FSnNYRDLmKTaZcbwjEaTyO4eJbQa0A5wy3BTPn8xz+4+BbWlyqXIt/R
4nAVWUBOUTnehXSxJV8DBlXEnX7fB7MGPn4Zd3hTr3n422//nea3zDyl0EaKHwOybMBUF/CU7reO
FoVLTYrbn0+uYN0zw29mQjuOmCic0GpgKQf934CoHtxzkJWLl8wjewSMhO/snP1CDAjfI0XHFhfM
KkBeWAlHit8wYY+tXXwQqnUeawBRTqvvRkZkcquhRuLqwY4m49GIABOii1uPztCUBNcbbvyVyGtj
JXAJvy6Rt8wgT5TKYmlWqwuB4f0lOLa45Zo9F+UVjOWh6ejtu6dXpqeUy6y2LFJnQZXE09ALfsWc
2YYE6fbmbDf9sMMq6XRqrITgZoni6u/LUjrvHuDlcG8mZ+PuDqjzTVf/wRd00hF3TMRij43r3Rfx
nFIF/DXWc7zHZsinchHT8+TbOL80vNWQAGV+2oW66SkbLJSBwdsbUpf3Adqns82SMJq5rE4sx+b9
P3dobtwKnOk1drth0ZzKEKShMzG1BNcZnyumzR4MwsR4lZD7gb7qL9FZ4xyRjNTaqsGYKLjYPKqy
egANn5A8HCImOyis4uy53k9gf24SB1xBL1QVHB3eQfg5N5VX0lASGyyZld0PSPxr3oE8dcdgtCY4
M5YQtrgqyE3bUJH11/zDNotFFU/ZqRbfyDD8gL2TamgIdlM7OVM+9XGp0Ga6MBkq7HdiYZlPWmNz
YgcXE07rPoDCFjrIx0q6S7BL9P9sw1fSEdaSv5n3jEnF+dVcXFxyRwcAkpnfxX0FxKd4P7H+aSsj
eDvO5/mEHhgjeAl1gIUgKq94qWwG74nzx1PcWDYqMX4M3gGG619BFa3GdS3iEHMGZyQHC7Qz7hlj
caEQ1EgqYOu7q9PQGqTo6gNqHLsxRftEIYbCtcsoSJ8eOlJzDF3E+txwzac/rYu9XJKVT+JsFKfW
ijr9gYJh5hh3c3VZQrj8Hc5RPV862/zFyqkdwf7GtOZzV3ZKpgacKA+53kKjUF/IBUwkI/vRwtUo
6Gm9taKJ0YrTu1bbQgHTg2aFLMuClAroziJl8AcjbQIK8gNRn3AeNGqtojlrmLYb2uhTEGdhIw+Y
bElpTb/bCbuxxxNqRoD3Uq4n/uEQNSCUxvAVXIYRbZM2bnowIqdF3j7urJHJ4VE+3TST5K/l6/Oi
vO738O1vDNfh3CN1fMOaYJUMIp/q2zgk4t8XiIJ9zgoj5m/agfhiVWKmdM5g4stouW8P/9gc8z4v
jWk2DI2Uh9mido5zTwvrkFtXPHVmYDMbti4UlYgJognJXwW+HCGJqLfcNs9cyYCZ7rQt2JWjVo1s
7BsbkBQCBdjgjq7ZAlk0DCjbDr9u7wy5VVzjywNlBvSltrowq8C1H9jSG55RRgV65DzrtJ2Meugv
JTTW9NB+7ObRedyUlTp2+Xmcuhwma9GzXpyKIaBk8QS9zE9WTE1qgExSBykn+pDQACo7z1GTHVcm
uux4MAp0pFLbax2bkl5gHJ7YVv+RbvNQvqpqTLPNxPRHnPyu15WwawTspPKa2/Z2Rytv6L0gsbz6
BzuXKTUUTZ/wCQmwx/xpIWlAGwr0iiaZYAYEbWI58kxdISG1OJAmQoZaLw9rutsXuIZAE7N2J0q0
chRhZ6+5g2hJW94PO8u3exhn9rT1ToqHvZwATtS0qH0Z9rvp8EAf1NOPk7XmnmzU/+piUi7Za2qF
rH5T7PwCpcPdxCliBGz/CJKYbwIkXCuI2VimwmNjMhQ2jOlY9q5VSyVu878fnVDGvx0u+gNJAS38
oeB9KSUWV4EEudynjlzEIU5lmEmMpaj7PMtCBLbecErDMHeB77MvtSmfEip0bPWIOYNd9vZzjx92
b801CoviOSIQpREVjoUNU00cdASA6fkrl4W1txGWWno9lOTgVKwNpChJp98YURelVC0UDA1tgZEE
qghvBjtba7Bu4nKYDNJBxwGuJpR38MwICDju5DSmirDWt7SeOixzIltUJ2Q6fKJK55MbR/c7l0jj
9fWMgJZbjfor2BR8qaeTwT38EtLjR5kJek6LJEY8UjHvWp+whSoiDDIplx4QmUJJ7oN/1e5U+21N
F3KZ40fnM5dqp1Hi8G0H+LSQKCV90xWeTIOHyOLQOQv3It5L5WHlAcsCayBCIkIFEOjroOh5YLuB
AhkB6gIdrcN41Hnp+nwIG65jrSel2QRhB8bQjhIufvZcAkdMZJMYNHlXBukRE5Vwqj28IO3E22/g
oGXFx4RhdMmDKXTV7t0HKdLyEjyyUg8pkYdUHiCMOz/BrvTX8MwQSinSEPIwuk8ThnTLpFO6uIex
rDAdySXZqSoeXGDuS4jMMAJ/81/2VJEDwKYbmDcfPQPL5lGnA++jrOktkuvFjYgRJPSVJmOwwDKH
43AdRitHJAcFwLJXpNo7ikNopQm51JOc7EYUyhns6qRrMmM2mkWNJop0miPRjZDhJMrJU4nh9pIE
4RF6T8NLWJhYmX+FAq/6MCv6VvcJtbbTSHWbKpnxaWbsbK37I4XO0tE5+aVo4XnHDHy2hrSiOqYH
a7m01VsZqK0Ez58Gppz1cET6rgYcibp7SP01AhNFUweGnH2+m9i/4A/L5o6wNQoOx8DsjBeTraMB
1OEVnzrw7bXJpG91JI9CkVMfihw2BFqd6KDv0KsGl7Q3LuuQBSMeZ5NMiFCeFX0eO98AVyjrM/rX
5fmp8XZUlc4z54fsJzNV6emUBuQ840so/6diTxsHWdwFpXl6e4frCerIW+b0gtTfhAu0oIve4qus
cOolxgH3E/ez9LhUIdR+kgG3/cfsjh/e+POz9USr3sN3vP8kB8jX8RF3bgPQkIaY76P08vhCMico
J37iFnLPe3qIKVJ2vuuYugu5C3urUudumvArM8tFVRuTruxIK/0cJ6Ss31rg/kimPvG/rF+UWHct
e4eI/tI0TTDC1QYWgsHLW1PJES0oO/h92XECYgI1cSircqQuOmzC/NHfCn7svmvHAUyd4na7BDmt
aMZgO3tpkbiQFXbAvCF9NsKFsrTUF33CstqpSoffXRgX3eUQaKIOEdzlMOjRr0YtHZ8QWAAndN0Y
pxqLkQSf5yHDEUpz9O+hnoAD/Pe34B9+feAziBRiVqWUpxGMCIG1JiYg01mNSE7RlKq/yTRTOHgu
1z8yAbCEi7og58L1IkAwqWbpVleA2c6m5QXxWW5HGTxmHDJ0njSeMe5GdVSFB5y/NdYdithkLUQn
QzAt/48f5A49r+S2bKwOhPrcUGAee+HODPSY8rxMcaUHqkoJHmNH+JN7O1LDjTl4+m3rz2q4JZCD
yrjUkvm+4E1l1JMtcrgUai+ufjmUa2mVRjW5B87TBw9curVhMGgJ5PZ46U8vcQKO1I1KI/rizjrJ
7EJxpMwCC6b9lXP8Rn+B9SgCZ0nbGfqKLhVAFRaGjKKf7kuWuDIoszMIVCVP5IKmHUD1OEat06WV
B+4soyJM8H0WA7AXdUYja+XN/+w0aL2qUJ0U0DwTIduFH5xocP3UUNaINg1qjJ10cI4sqpL75515
DUdn+5V4lFcibF0YlsDgdtNXKfUtG9FRKCSpAtvVARki2nb4be4T+QSP39idjg1cNNOVdnd0KU28
f8+mQ4t/NR06l3tg3t+WDn8CYJ8kJHKYx+OOULfBwSiJmHXc0d3b2aJ5Nuj4r39PLScSzVJWbevN
Rh3aZvzYNJBH4TKn9/oYv9eYtZQ0nkxsBHU9j0Ope8/rGHAX/Xvkb6tvagXnJu1FOOFtVhETl4Sv
X8yYOGHIgAP+iL5L1XbjyMpcMvneSYARJn/Rtd3SptmL3a0GYC9G4QRaG4rDpLqtz1WRrjfj6/qm
zrJIB9FwpCsSx3Y75lrWx+nfrZhmCNq3yHJkwO7z4Rmz9xwE0a7/R4SZ3CJh2l94+MWgQc8YUsTS
sKrIJqc0ar/pTMt6bBtyrxYw0HXox1RbW9cmYXp+947gGdLYBTo3EWGzkJdbaj1ijR9pAgYsHDg7
wsD4eOeCIJVBcQPVUMJsyO7U8JbwpJiyaxPcVPtGDvznk+vvH1S/2G++Qu9oeor2raNlDYBoTN0a
L3onxvti+vxMzWyrPMg5THjtx+cH+1jE1tLiMHepFRTxsne2IgQVKHPpQX6oRx6B5p2OJXzSpYde
d7i1wTLLYbhVs5anMXRicbMwckdRw7OdL7kiBZFt5cKJUAG2KlO2O+hBgbTVmuV7B/Pv//ylf/F0
rWD5TxF/8F4pPkFDlpzbxiAjesElp8xUFFYknQ/tMgCwyeGtlzIB5qU/8ygT943RZktwwPTJMAko
Hl4j+gWrG4orRzx/8Ifm7iBaHgJfdncYEIiQOm7ck8jr0xxRYaE2fNAQtsKX54R7yySgCH5GRBj+
fh+PCQZfz2iP4Xjr822OJsFIxs3zVW13k9OsoLNwWxCij1eIsWnzFIANUfYF9wp9q5HUDmTpT0Jk
4pmoNatLFoepjSWY2mv63o8TMn3+BeckmzhuubZSEfP0un8IOviD2Ho7MdRt92IXt62s+VitRZaH
bWiMcks9wMiBlNbZY/KNL9PfaUOFbo2GYpqo5NojVNn/ONT/oM3FRCwymXS61FrhCltnFghuiI6h
cOToQkxyqgLv8zXYLeGFV9hQ+k+rhNjXApwNmMBey1nJX/F5X9qir4y/twiZWn5hMsn5Goi7+78B
hKdC0Q0mprHkmq9LSpyXTDcE5fOXwPPzV8HPlahwW8RTk1Uw9xderNrSoBdfdz8zutDn7Iq6K6j4
bLYVUWJ246yzOWaJXsRuhHQX02uzc+pQgUlWHgXrxDcDyWS7sYOL3MwbGQadgo7S3WQquEq2ILXa
jIEMo+ETjE9EYV2MEmGpxMHkjcSa+WqYDDos75B6JpD+PAdAr00Mikios3/kgN9VeAlidyF/2Xxa
/qLNZcxvyB6SJc9bZNXlZiTW2JL81DRM4jXsoo/HdV4aICf8aysSYito0/qY1GLT3TXEIn3By3GN
QRZnROTxi3Go3XyzSmKg39YcCSH+Ktv3lvoXBXEECUA96C6yC+KXZOOzIf/iR0B+j0SwDnbfFpFY
TJtiF4g3TI2s1aSMVSsrI9MQg7Yd4H5+r0Dn2a2QElWdhjXIfwNqUN4lLAXiIgCa1rK5tte6Zdld
uCIuNZhZxS5AB6eAJItwSyA1DdtiS/hz0/K8PPDUKISxTiJf27sZY8Ew0RqjGCPYyn7FpxsmEOjk
YV6BlgG7TXHQ+vnH7Wu8MVbMdU9faSCSTsqR9ELthARe5BT2WvhwEu8Sjh+/98xhou36hgnfdcTb
Ml+2qIqp7+nKKdIgH5FiB9PyfS2JloqcJhqheHb2v1R1B1dSemfeA2PAw2uP6fRviS4eZRYoW3f2
cSCBCuuo6v9zEtVVdgTbUoS37Jty8LmDjXJQJfgySqWpW3wl7W5djfl4X7VI4gU4UY/KtRANSUCj
J+n9tUueZNwd7eRngNQHzE+Cfh4zdlOI62afxwN0gmrQBWMtFxdYwgy8GNNJJ012qQBuujHP/ST9
NJkD8X9X/4oNMNa2ueJDW2DYWVkgqjZCqxH9rE2LSJwiI1MqyCPGkUTtvgF/yyyMROtesQDBkjWl
y/W1dF/Vx9iijg/6+VlxUxAH6335/McNyvL6gBOVVPwnUdYeu7nvu4cnLKP8+B9AwcCb0vz/bGTS
Hl1SwpaRx+NS1q2S73XypA+8tPVhZomrlky4V72/UkEAcd7QSgaAAuSd7N7Q6JbhX2gp4luMGj2o
B93dGs48wJ5nIvwq9uCpLtWxMHbNUshvI0TKVD/GD7uG0CSJ650AvoivJ401oQpphewt7lgrCWK7
1d5/P9BUM45W5raYLoIC5VN///FKfHtmeWIx8ZI756e1G51FjIS1WuKgoKBIvTAyJJO8OKt7H0K1
tBn5VmlK77Oqs1ogCYD5JEiR1FRJvYru9N3BpuZIrxGDJ1OislKWtUqW5v3u+yUI82pzK8tm09kv
y/nMdgysZ0d1njbhK35tJEq6nC5RZN8PmPZZQQL3QrRRJzQAs2z4wt1pgr1WgHWHlOwseVvLU9/g
a1NJ3XteU7QJ8y/9z/ivj2uAAHj7iKAZ+hBmyRQaU+StdPghxu/0wlYCt5D0K0OBFIvizfpTzcY3
InMNibvZd03swOt3swedJHhwupRytO50hRm6XvqCUEn4JpydXFW0XMA9e9VKVmL7Thv3dlZ2RZe5
2GFsWxe2J6VJO3eTC5QUnuq4ARHqj1GWpoeoOK7CNj848J6EhFULD/Biag5x0/9PjFrSRAG5hVKm
s01UEtZN7IqNAptwrSO3QPzewllxirU8ByMLzY62CntdUP0HxxbIbgsjLqFRgopXi0PrEfhZUhDX
lrYWLyjPlZGscMtyDJ9F6JZ7BU/fvISi3EueZGi2NbnFHcQMPqFfIdkvEKNZMqnt8Nfp95yWV9nf
tuoO6XInPfMJUn4f+i14elo+qGjLAnalL1cZfctAkkn6e0cr6YQNImJBGHuk6s3LpcJDowRecJRO
Fd2z6OMflhTvCyE+64rpwet199ihD76kYLpZkwPnxZNmegoHhnUx6Yzna//SJ4m33xHIZgPR//0r
FeBCeJsnfHqcEx/apT7ua29GgDsTkG4oKi+K+404jxfew6ExKdeamHx+19sAMjPr4CtcjaewR/Gn
Qd70RcLeZ0UcTGFAdieN1pLxESQrQ2dKoHh2VVgILX1LH5HSNn1YyY77Y+cBR5nDbIARQWMWSYM9
bgwWnDczaDA09TubjAbEHm/wuA0ZCp/KhqAx2Dvduf+ll+PFpjegSTrUTEXx/gWWgyluEzjeucie
tJZrmcgigWwjAA2EWx1Mpb2jXPf+5IVd+/0UjTjyia0ZRQKjRPKR2bRVZL7kcQ9kEWIXjvJ9H/9e
gbQvuJJ7dLpUxwKq3RDWtRz1Eq4wkRHIOy+32i3yLZeZ56fjDOZ/2+8kESaHiBqwQkWkw3NdET3C
HzGDGDb6v9q0vP/g8CmCTL7u2T04xiHWI7f+Qg7wZO4FTOhG71HYq0Jhst3aIDF0ct4rRfLubu5h
hSpkEVJCQruK0o4IGavi7wR7dabpb3NhOmBjmMcxQUnOQpwcGJSUh1saNn8oZTozrer6vamr+Qdi
HqFAEejMH087UnEBNYULCzkMaq02zswtswzvjyCn+i1SI4YTSOKBf02CILWUa9zL1Wuuws6r+p+S
eWBYCDXib43+UBzH6TfHmPGrS9w+V8Rc5MPztTS4JnMJpNlx+uwk2kEPeEc9VIMJsbh3pYrNEMR1
KHI65nze81FDj1GaX01bVA1aaE4aTVeKIzd3iuhgUSfkUt8/npn2J6D5ljYiO64m6g1UrFh2Odpf
aMI/je3n4xvA+D+dAEHpfa2f7MzR0+DPKKJKEYR+KXG0g8IO7AMOOtV0EBVRVRopS5rKvts3RdMh
4B5RVJ069Yy38288gvMRNWhKMdTU4dkFvlvB5rjG0hqmHWFmj2wozLzcnrYTiwB5It6s4WEAYye7
V6A8YikovNbkLhKPtSrruQ/EFjiC2XXskYAdyfSa2t5D0/IjzeFhJhc3QDIvgkG3YWD6nA30Q0jR
Q6KOX2OJA7XO78gzctw/ZYtHWSl18iVF0MkNvTqhU/oSv6VpGfQbqZeWYs/n/LQxGHGk6H3sugmw
JMenNrlblfzRoPcxUjQrXdjsLl1ohkMeLAX3DSMMb7PJ4Z2BB3EOuSn6rRuFHudUIx6iwg4vKLAo
mFNlbMOgLVuWfnNyNLYiQR/S3iX9iX4IPRsDk1XNf61QRaQnmy71dfIt4AI+gjHWaQerLUTpgeWt
1AgUxUpjp+aF6zgeMDaVS4SUBuSTgNFiJfsqYGAy/s9RSnqtl8hh2SMbEYB1BRa0Sf8RUvamMcxR
KNSO24VAxS7dwgxUFGvbjaGkrxJlme7RVUCQps7nKS93HTXiBg/l1n3rI1RL0AWYTP+Dx5wqOhzu
OCBp6TD1hWdK3h8zPzuKz46adAShtJdkwcnhxcHhha7rBvFkigZhEmbQaS9D7tIOMGHbzgc3Igel
bLFiVFPAODjMANkNohoG54BR5VoGdGJKgCpEtdobWNar0OTaE0eyqe7Mxmb2bGM2bSn8beY0Y1qY
04WLWJVNbHI31ycWiiULiVEysIe2Qemr9Ov7aoSl48ydzBQs+XKC5t5eHAzbcf06C0WYke8SCJTz
mw5CkyRGrak+WlU9oSQ2399MotRmeCqHA0veGKg7MI7vg9YDizh89NiOeGOQ6nUQ1l9DNGWfKtnC
cVyLHrXusst505IPt/5K777QKaQGv93b1Ba1StShkS2dMYAJf+SOcA/RiNAj7RJrd4jL6WJ5DoKf
CMtNrGqHbCOa+TXR+Ke6Vsj7rvhDMYvfNP4+hqSdQRl9B3NK4BSCC6/0S407BFhlILRvl8mOuFiy
vSNpkCG+9PZxXgYvV5nvjHkIlOg4oFrafVYDziKpkXrDP6D520wmelasWfAk6wIfqu/GlERQZ3N3
/bNAeoBT1V83P1WIR9+058tKwrcLUQS0wuqxC+N9gcVnP4MMN13s3esRy71TzNbkMzhQNtr5IB99
QPJBTxnve034dNV8Qn9tx/iziTyGrwH8AkJW0GqZUCECviLjc0r0PPcIuUcDDf/Z+J2+FNdSLVnr
EDL60XuIE1H14vUT43An9rltU0i1rTO3t4XXpyTCWPip3MFI3hFSR2ebF4lXxtmS0+F7PN8w2CAO
90rmEbBB5zjahd4gqyE5VBTGHRUPmWWVMihyQ8KpAkg6AmWA3wj8nXfFAZKEF+CkUcZu7jWE6KC+
Vq1nXzaD9PrUGQMVVbQHN8iA8bUR6zvtKb3iVOzisQGDVBi5yNSud1L4a4zTtiuPijYs44xLR8Ik
1J31bbziLDE/M19YcstbtLNkV/8Cx58ZwXVcUcasxBHCGHb7tnySROz4WVn+z+c3Eyv3LFE+QbKH
kfoewhkmeTtQMdlaBJ/ZYgoMXPGEFoq3x9rgIMRar1jI9FbFkLrjiV+kXqHabkrzrIkmhaqC4FoA
4hJ22YP0PoDi0QhmY3hLTamYhUXvR3KfQMNtGiKAjyJAfK31Tfl/3lJzyOTzZy0mGyCwgDHp16AY
YY7ihgk74yK7Gg44sj9LRXDnC8ZAuendSWHLbnCzZY1BnmF+pIGAQ8HjcPYWw7A+dRg0ictr/fDQ
UVzP0f9XZoLrTUZHn/XwYgVwzUilRy2awl/ExyqTOSalyMh77TiwPO1z59w/3mt0RkZtno5uGi3h
DmuyenRGIEyy1N6fOYLrezYaCeH+ziMT9T5nt+BirFhNWVZTB0DC+xXsGBUaQkdHvhb8igkzYuTz
Apktu9mAaaTqSWDXdmVchBswcehiXh0S0guT7BF/1cgZfyT6c6mjsgQVzljMU8j59hqLfzoc1pc0
2flFJj+igAZw/MDEHtDck+tvfVyz/OHZXYiYjXYMp/njE59/Hi2Y9E3Il13e/5MasZJH26wOnp0K
2eluxcgDSNoGvbKehNDOW6sJPvnGZB+JGG/wo0ZlQHK0UIi8Vp9BFrGBxiLf51vfNjyP2ZtrltFA
YlRGRXwuTUp0QBVncUoZBzszFcDuQt1tntX5loHCfD8NKw7XY9FQRBI5smJYjGFtUF39VhPDHzAt
CkEQKVDGCZvOFsZTwdwoHtSR2/ErlgqN01wYMgdfTmL/zBW/n2kFzIGSJrW3t6+MeWBRBbRQArQk
FVRyu22bDEq4+KdO9qGXw+rKMNnYx8jAkIuaTGWANbvt5oTwCDegt4Z0Iz2TW8pSfojaWmO3GOEy
sMYzmGZIzJ0aWEtz40ABF7lbvbHp+xVBX4SpcBdwvLmr1zBHVKhK1mrW9e3lmdF3I1x6vqEFh39m
sf2X9WqTUhMQfLtA/2vEBwi5by5+addTSKUYSsogaxtNao0QYT1wRnR/MfsmImDDJJRohG28vypK
oWO1r6C8qd1fV3ZNn/7IaAHbcETijDsJidJHCWjNkZrm4uTHFYx85GH7yN0wFkc+nUe9RkTG7hAU
Ls1s9BKquQiSGctwee2drxJ+gwQG/V7nlZ0hIYMHQ7lfVU7mmYzozUEKgqqzi8VT5YjvCM82lbC8
g3TRpXO3aIbS3vXdAbjcZgraiwlBhwWwMAj5S8ngCLz1rOSq0vqitfouSUdDixRlIWmwCDmzrTs7
LtT+9hNdFN66ZeCnIwn23feklPXfTJqeYRSgM/yp+s4VkAa99MjC65iwI41uPOUcm5XmZzQfN+49
5Vc1uDWug7laoYD956+mbof3+I/tzVcCqOjT4ugoqK1cDTiwORVJR4u9/7sDBGtAYkYNwXciqD36
BKiqxAPg7kL1btFGg9Vc9sX8fzxiI+WcoZnpPF4GxhP7vGHJD8dS/LB/1OKSR1tg0qyuraFdtYk0
LUmN0jr356J5VeCQTs5V+EMAii6x0+d5WM4cYTq+csBTJGUbhMzo8PiMT54/T1Fb3RzkfdIp30zj
QYuZOuRZ1lr1fYhQCW6QReXemAkWdGDyP4YL8MMxkL9PrukHL+s/Q7O2nLuqWImj7T/PjwKupBNw
wJlTs1X9i6mCqYAw88EcSHXMcZWGeOmsuyVFiQvF4qgzCa0D7D13Bs2ram1FlrBmWIKBFy4sDZSZ
YAgCkiZ+vFqad1pnz02Af5A08IhxZLGvOHLHix8JL3hblRmULVcdAYHphCxapr7Jbwmymro5ot9P
rpqMnbZD+RXr+W8ik3T9mtB7iGUJXa3eHutfnOxzxAxYbtiIWoaN4P+tY87c3IZhm03DZ/j3GIQ4
ohkH7CppaqWl4gU458m3P1iBx/JnUHqlNQx61Rr+MpEhLlNkjhvfvlYtCuw6yXfOmcWAMs937vqS
5FdjT90xqYqv8FhlqsDo/lfPj2J5X6/mAG2yFYVwd+/J94D8qBu0s2TShdr+rDec+3E/Orom9ktW
5PcLgj8M0eZB6zC8DqXg3zqB50ceGt1dQ0r8Hfet+nsl9OZkx8rZbecw957gGiM8kwHJ1zudJmpq
VW5ai3CnrmDZ3LXmQr2vOaisUvFOXMLppCJ/cQ3MXbGe8jedM7uOBJZx8zXbGFseDy0J6itSfr9j
6MXK9967BeC+6EVs01uszFE/FZcOVqRQ48DdQ3crdFa/bl4geo7JXT+z3x/UnZruqG+ocsUnheF8
xjD2vHNANkPTY6YtBjBCdQSZ2ErSBTee0jVmHTOVZR7l1Ha5aoAYWLeNbttNCBt53A5vERQTb8ax
MeY0Kfaee1/AqV/1dR7oIuCMaqNkRfz1i9ponp+/sLwi5SJtqHH3Pz1jF8IntF4XRyQRUOy2m8P3
ZYg+e3nnwW3obTYZ+M0UnFeL9bMU3ylPAXJrg+ZlqcwynXE2kTlVJ7KAuf9zvGbV70CpYIBS/t6P
Ooa20kuEjh5oFewkIfU+zWo8gTk0zQeKK/Tt8ZjBjYqqh05HIiFM7IOau4+ZBRmEmyf/fZvbgimX
yAuAwoqwJRGktVI+VBObS5OITuu716O7rB4L+7BGoBNmD7ILFK6A3Ksf+JWFw/PpO0ocLHY8H8gN
HOrH6ZUGGVN8DpG4aTRKTlgPWEU8e7kCEQWQGyYme3gLV+FbI1xS97vHe+iBLDzTOFC80NG+dE1t
xLNj2TGSMYyy2O8sOaQ+tMkSc1UqPB68NMk9DGSCE7DCUSd0AAxeK7Osmj27xI6JhCnfuYmiD9LC
WK1yoXtehMwu909+/3iyihK0pb5BxQPG2eN8HJnOl9uw/bjEOmHaVSTo1IbxV1cppucg0AZW/d9e
ORYyV5mgyMfqggMdte6gVixhYvqOgQXdcIwNf6ml9krm1myO4O7Nyr1iB/2e2crwuthPQnTMV/Du
853WjAZVQJ9VON5dLHk6h/auWAf08L3llui5K6JF25zbXzSLq+jo/+XaMQCM6+eDPLeeGb6xUINX
w6MlBK1uYXfEaUIu6kFhlyzuBPgHjPUj+aPAZ11Jcpw3zwlMGava2f9oq8BUV41LlmqcRzbZu/UJ
XYKCxDzpiVDIljZ/21Vj2/Sah24Kce8sUNuM8NbeIspHTcchkuz3G84jCYm762jIcZhgmmShwynP
IkHaD/AnylI6Fz/x8yJc/SmGLwyI3OK99fG1olvKAFReHLeNiJZ3Xjat/po3zfuE03WQUYWbnq9F
tC6KvpxCfOuPk97nhgAwHjcHhvJ3LyfZlsnwlL6jUs8amQ1hksI+Gdsxod1amoG0ZQZygpGzS1cn
Wrnyo73Mjpfdsm90brv8VzP8frIIJLgiihnSq5q5govdvxCs0GWu97uYe5owi20aZk8a+Gl7Q6hK
HoPI4eJy1K6/D8PCimmwrmWGWH4O+8SozjYb6ajNM1SzxvEv9NMRicjte9VcKgencdotc6OXHF7F
u8qwF7FZB2TmU+yopLWkJE1hnRQWkjZyGJSdcO1h9RUsQar05yeDyvZ3Pzws/aK/t1DNnsDZNt/D
0AiE/XvlS8B0w8i/UJOeK54VFpzxdhclL6rJ67cWe4kGr9uULfjP4z7gp0wW6o+5DlFH/HGAHdvW
+IkrTZiL0BYFYpcpydhyJOmvaYfj9oezNh9spc+CsG17x99cClcgLUAYSEn83Vz5ACbXrOqYS0K0
tqzaN+/LudjaW8TywBsQcOz4pE/nF4PWvNzhY+xYD11Ip70vrQwhgyIW3Z8dQ9fBgZxl9NkxacmV
oWdmmHXVcfVSq2u51FAM1E07CWIuVQOozDfucaFcbIVFy7AB4ZnQMf3cDBMhSkheck8jXC+0ijus
3/hzg0s1BWQw1DXI9+Kkob5IRMeIDlneebgmiBd5S6rD7b3N9EYC4GFAltRpU6koYDFPGKPiXzNm
z7VsIHEnbTYfxqCE23koJIj6qtDkF4GlhaBmrPSsyNwBw4dFHs119LTamu1ZuVZ7O9VKgUxi2+JZ
GwmPXKEocEve9+Hw+QDl7IIuTKhOmWGTv9pT25uDYrXSMxBVDrpDB/odsJrC7oexw4Pw+OnkiY/j
d05loeKL5sK2dZUA6R0n1asYXLp3hyKi4QdmCFHJbf0T3zSOnsseyTbNQfE5IniiO2xM4REdIQXE
RjUJZsIxuqkH7V0yPG154kDOMfooCTBo7oqODicNVACoT3Deal60cPnh9ta0D8RjDtelTcxK4PKf
3myXmjptvpztBsd4DH6HCXkXuoAV6lwkrdaPmPW+1PdAmPJfT25X76SLv7yWduWUJcozCnHyugd4
m2gqVGYs0w0xOWM9th6iTZOmHMxE17bvk8LcyQCcZF+4WDfhf8aKsxPqcus5MCU4RBqdEY2J8619
BqILGd2FHpv8O1FwWJi6zUhskLeAVmY4Ga9i+lPEbEvOIpiUxJQV4aJdhdT3HaW8o9JaGYLx7riN
l8rqTRLuWIX0oRj2e2F5S5FWgQSv6PH3GNm3Jy69nTu9rZefZ1/ynoycXucGvYbXKStvjwnJJPhd
PddPaQaZPUvuqXTFvhrX7r4edAoFR+cbORUz6WCpWM8sLAp8+59Dse2bJ3heFqjzA+OC61YB8oPx
MUOhhscH7pzGO+oBMAvJfDDoFmINPk4y8vccQouIHN1bc1OSW6jljSQGPDuZn7cqB96e9zwOZIJm
MtNE4f+Ga29Uh/RCFedglPENAZerETfrvTEtyvmQXJ/nsdMEiD0Df9VKsI9/owWeIElgN5hdubdt
YZqC8rlaoMBTPsQzbJfvvUMMbyrvjZmPP/0OwZBEuPm+sWh42dT238ekgsw+8ZM8b7jSgb/3gUGH
jIHjBgfiPjBfScOjtylgyHkUVzfLrXf8KPoGI1nfDK8JesQnY988D3tMB/8tOI+rvPGM90aJ3bEM
71XWZy3AxhEuNQF0sLBGIqJCt4JnPHcEbGkxHJtUwjORvsoThnbbXUoyIIzbx11nZu8IUcaoyDgm
wSAhd+O/COxvCdjc2qkCTilZIWagukX+PJFFI34MsmI4iuS3kpIaSITtXX/0FK/paLVCrc3bsgyf
Y17RZQ+TbXw+x3Hj8pqCuiPP4FyzQi8xpXVZcpVb41HETxmbvlKJrkqxsRt1/Isxswz0w7Z9V/mF
NpgzE21vYBbCe64VIkO5iSaHIqxLIeOZpGaDzWpkBmyGxM3xf+FsGyN1WckN05EuI3Upq0ZNL43r
hKK0G2ouxCnOifwE1vNp6w99Zxi6NNynhLrAvupc9RDcc7th2+Axu53FaiU0DuEJ6an1pcjOObBs
aEsUT3c3fwKCBtPos51YySQAUXN/fCL5bcuLkBpe4buDFFSL5m+rwYTt37+eudAZKqz6JT9fbw7n
EvXU/0pmOS3scaBa3kdOfDX+LJq3ka63xfvJT9uX2HLbYh1vmNUVYIjr544snolPtlJdK4X3bnpY
Ic0gjBX61i/EX4JPu1De0gx4ZMaxhjH7hg9EbDy2rDbryJi3szn5xsUSpsK5RZJJJfjBBRvjeVwB
xD1ULyduYoCPrEXK/AlTfQ7d9YH4yjdhTULmRHdzE30lVcrQgazNWzZ6vmWx0Sk2xAYOT32rP5kV
VQbZXcUxFcjhmcWqq1j/8iTCCzWX7QiJp9uzVbxsV0N/v3dMtnOGVI70HcnDJbeSzThTPbK8Cd6M
KindaHbwU5B+zpPnUf554RjfNeLb+Li1cH1nE8BCKBa57FYcp5jE7IolKtAKr7r1bNHhhqPuVsre
k4WRbEG7Hg/0GFlgWvjWS6VCz6x7NoFM7JRWcQkVo2MpjKybkNhO694Bc4B0QwezpMoGAY3USBdC
AGqeL0MJO0djHfb610Ed+2I/VmdHMQJFwbDqZTrTRZtq0hsTvwaG8lV6jMzq8D8G2nw6EnerEWZu
eC7KEWLeuu3dy3wEMiftlJrWu+FlSgTSIky76/BB0h/jvKE87CaFTFabri55FFvRM7wQ/0fS8Xrv
UMvERJvdy31B3xTDSlX43iTQq8bUEK8thqRC8Jwy1VaqA/8Ym4n9b/rDAGW3ExHq3S3f/rHTqN8W
Ub/Kvym8Q72XIqZG9jUIw7M/ihXFl4d3biGLoMzGPRu3ZxwlAIXUdK3A5FYdfsAunKgMRzmLBxQ+
cK5lZMNmpOE+JtGfp4ZtGQhpS5UECCFoK4UDYFRgPO2CEwR/1qLJ56Fw88+o9JeZfMHSsR4c+1oD
//ytBZSfoLVJzplyUXmBQbQx+iRDXPIktzpsnAItb04NRWIBmZSX+vzAFBX3BToJDv6ymwJ5Uuqe
LaswEB6gDDgt1J+H7eIbxZa9vJN2dSc/pcJwIh61k64uT3bvb/l+C9DhAyQ1NqTTqCV+rXv1Qgij
WJF+dmT9g/YFnHxkIbgpT86qylViFtsLulXa6eI20PFZa2I/xNsJC7M5ITnA+imUpU2TXukx8ZA4
n419I+37Furr0MzcFZB5wq3r+I1AQWCX8XYepBfGo+8FVHz8SWj4zy9xynICrz5JG7yWFaYuRhl0
vUrX+N1kRhmaQqI96ueiyA0yUSDVyPuM+7nyruKXcjaxbjJFFO+5VjQFJBZyAHuqc+SRmb7FbByw
S7NOcc+KLmoXHgffLofwOhpYn+bnlcB0R3AcJR1+Dh88as2/Cy7seUYwjBnTecB/FyRzhzW5I0Zd
HLFizDE5/M5GGPHEYw+kGCSbqs1JcKZyiE3iAU86F6lFaSvn+dz8Houa7xqCOycN9QY5QZkFfcsp
Fh+dfvQsqszvM3O7fPrBHys/m4eiEbbkGZMRJvWVUaMuI1m+6sBApDCX3UvFS8HCr3kxVniCVe4m
KialZzDWXxmHGxAuO4tS34xwdIo4MvVl9mEakOfepbddcBDG3VXfz/Gwp+IGgOlvroQQNLMNZIr9
D/vPNQwiLDtsTO58DllyjMM6qzgYmQsMY/PTVGISzShMC0d7crgC71vGkaI1PMJuu2Ocg60zS18a
fwAiFELYjiMixKXd0aMDN+jZXbybsA8f7MkRmT48AdAk3TOj3ayW8m3H4GzOD4w85WuhLw2rA5Hn
2XHB0Ffm5KjfKv66hy/HZOT58sudFi/eNWAQa/OEnsnrBsx5cRanr4zw6fyphrqcJVQuHOGj7IJt
gchQCrLlrILwIKvKXx+c//OJFfkwiJv1+HwQr+gYDEwdvqHNklgbFysW9YSyrYAzjuCMfc44O8qf
gjZgiex2mUy3FWqQWoK7Pzemh/kgSl6JgR02U9iQ1jScje9VZA/T42Sg2sRC5k564VxOV7RhNClu
4BGd5lzpl9aspjmu6alVel4+CUEJ9Mrx/VMtM4yRwqQaR0/GuhSZUnDcAlbVR5rR5G6tVC2gtDzk
eMURGnJeD+PJ85EBV3No0eqRLf1nCHxraXbydhh1RJK3vSUIR4TRVn1jKMM9VRhqr/iI1XEmtl55
q06GgCABp5RGvuwp3jmULPNtrL5qNmZ0LcurLg4zFLpCrvx3L/6hDjb7poelh/kWnOyqxJw98g6x
XMNIP1S8xFpJXfMxTDbdNeOR6xE77Z8vZXrs3Obfd1W1fp2+w9o9sTVAQbVEaMPP/Of9ZPIKncsA
oUs62zoppc/Gw7dZsVOQrGxVK09DjN4GM1s7ZGTpqsxm5l8GeJ9iG6CeNlJtfGgj+T8Pnd2hrj9i
XvL5QR6/sIQ4Ld55BGDd8AaB+XMuC3be1RPYpWG8KTS/rAsTYWXgvJKwbkDRzkiez9ItUXRctSu3
EqIhz/A8HobotHKbrZR6FRDaHiDu8bHFostgPa++iy3c4UlnAhxE1LyVqyGvrBmuURua7KXU9KJX
3Z1VooBw0lEY0pN+M32KygmKOHDLPS5Qv4cwpYIqC7Zho+3K7FPEKKdyuIWjMLxYvV52+/eY8NOu
A6/6t06D80/EsdFWu/v0WSOnyCGDctdLYT+34penAaRrXyCWzcDkQn7I6rGsvfJii/tV8eDoEZaa
IZJHCZlsBGAnE8bsaRIU/YWtKOls3pcAI6Te5aljXYHDeSJohcseOgmi6efWIbkrgXaDvxzcRK6f
79hqB+FDo0VXFo3h8okQgfk2yoTZkD/Bq7liUgf61xazU1NuENTsQKDtfPP8xi6hxKvXPpAcklTK
b0KsukTfVd7vpYdmiU+ZvQTB4LLr4hjDkH13n5Epiw5Y3VL7dA8jaqc9Fpq6e/+JUAPjC7nu5qDG
WBRehqsZ2Rv3Y04UQbQYgLl5orNymky5cbdaCe8ICZuImgt3gSMiqGZfvITZL4vDeVsqRjh/Ek/r
U1zoueOmQIf28b1txQ5dCkTcoADgzATTIE9OhxJuNLdtgA+Fj4SsXAIotD8I1pIVdsf8h/ij0ZWz
0mGnn53dfS83P1yAJa4OBHc4f3iiqz4rZ7T/5/MKZ+seeBo0xXSyImCx1uz+9o7LmQ26tuvcgGLD
1ETF79APaWLcFHWJAGp4AtctBOq6WrO3bXijv1H48AYTkp/dN8DTaLqCRCBNMCe6RDcFUlBQYJFq
alL0rpOmOpNSSMxwUhkEX5vdOz10AHFmvE3dLUJSq/kZKSOyUgbdoEwGRGL+IsyovI1OQOn7gtcq
88STSeHcnfh35eUkXVIJyLNz0PXDIwfYl1+Nst2kwbNmHB9aXwFG3vvInYb2aM4no9H93Q2HABMD
859Ne8lMCO0ZGHUSTV6Dgy+69bQ+fs/R2E/UIDMUeNJaBlt2Q01+nBTVHZKNyjoCn3pTJ7XHy/K/
PFXLx44oPiYgqmLJDNAyhTu41c5TuL4ijdS2DpzC6PrRbR2Gn8HNC3KX0z+Q8OI5Ps26WyceL1O9
mRMNngYAMFlx7lFrRZnEciLz4H6jh8f+ax9e58tH+t3Tq2o98plUok04VwYTRenN768aSk8R+AbZ
EFbXY1xwSEyQ5sbUvgsjGjmux62h+xEdp4FW6DyU6wC7p18bCLBbWgV22yjU5qS1ggLqgzWa4/mh
IR5crbQZRMlOku/+5t4/embNv+y8Qp9ray/tWA1y58hL8BCqy7g07rssm7cDzWwsbWsux5EF8i4y
ngn3v9+GIQEgEK369zCG2G0L/7VjyFUmnLdvEvKnaqKLah4RIn3gfWV7obGdpk/wm7Ew5fzLdiRV
oHHsb+N8WbzvXM0Y1+ioSW91d5I74s3x1Sxu0rEiI83Iko1KfD+lJFr73izjMoist0PsR8IkSvr6
z4Rup2PcWrUahz5b6WgSc09DcUsYYiwjgEPzbW7Fsusy22QoyGCIegyPZCrP8V5ObVfztimSxvMm
MEJpen0Prqfsvix28rBkfSeI5TPJVBffmsCn6KqhQ0k3wX2FKcSYG9bK7HBTfzWLpWhq1elc4nHd
vEwQQ+SONys8egSrMwBgKA2KmqIRbFNdGoxZBYbwUGnzipwBH7RKNb0dOMf5KCPNYPw/O7RBUm9l
294+Q7oBNMnIYF7T4h9JyaCAbbr9eDkS1EjI7DjGPC8F407Sdi4GdDJBV9Z4mv/usshxkL6bHzba
CRp7Cb9lsR+D/bwqC7trgbSYN0Iq2/x9olcP9slr0sU24vXY+U8eXe4++hJgVqjwMkxfCe0OcSGQ
nT8NXXdW1x2WEJIj3PrsSemBLnURiqYN4CZ7iIaonhWM39MNYaZS6R78MdIXjm97olux2aiosdZp
1AICL7jA5UqZeXruriXtQe1u5LHutwauttXu0+Rbch5vpdLRVOyXw0uVR9UBHxbuH6BGX8kiGTXy
V7gz0uEfCN4DNMrZbIqG/StkGN7royYzVh1UdjjmiHZ7RxaUISv9WgTf/GcIFKpTDpO7MWvJWgv2
hzONG5yZfKHqJKAn2w+VZe7tjdouo60NzuffCWRX12bL/jF9PnG4QdTY9qBpqTHpVSzIWQV8yUy+
fMFDpwQbdi/kZJ30oYi6CpZ+z5G/YXib87rVuH4u67+EiHPl/XmfFTbaTqF5l/DCy36oGgWq+US/
b6X5iH5EZnuGljBEwqfnxmKtN3yuy8coOE3/LgYyuqR281l2Nl7xXFjP6ieAIQ3u4gnaOpbqFwuy
SeJzyDTcfE84nKcHDk/JW3fVZCzE7A/85DiEyTUgnNoyegT3GVkyfNxRuCCupmOz3HLUynJ+Qvkh
KUGkSNdau8+r6rV8dO22yp/z4A6p0Uq1h69Bms48Mmz8/DgqRSSjSN8TKB8BTs6sONpYhPa9kEeo
Vtam2gEk9ZPWVQCvjEJitgEzZsVLKVOV4d4qywAPoZUVmLUGYf39Je9Kc+MskD0CIQQZ83nOlt+B
SAczjpbo38JJQzTNFvoGcUfWvL+ppiMvwoRQoUsOvBF1lnDfap/d/az1qn6kqXhXF8WAbsEibu8h
c2fuVQM5eZ0q3Jk0YqTOHmkVPRubtUT1+svt2rGq3NoBUfWGmroeBC5kPQoxm7BNTI1wW+ijhYry
y9Lp3t45+UvjQUNvJ3ZIY1B9Wrn2Dw3ofGugresTkuuNi7skkonvaTfStmWrnVllG2C4cLntxH9I
+AxQdTV4nh1lQNZkLxB/3aStBUn50Ky5R3AGDfQ4DPWJUqA/ZGUuIIRkfafHVcv4DuRBcl9bx+Tb
thDhqpcImxCwzy+uKuc/EjxevA6azN6L0prUHYCpZUKt0cmf1p6IYZ4nz9fvkckY6w8Zll+KOSgg
QVoyhWUEYwexhzQhLFCLsGNWPKgaeXFB2Yw2+hiTwp/dKTUnbXMjgCrLYXSXKqUaJa7mkwf19iEp
bKc3XLKLb1ItGERtKTmTqM8qw1gSOSdcLZ3cb2DtmXVg+JGz/cDevBBWJ5FwqqJErZ2VYWzkP893
QqFTdJZKzxaK/v0N71ahZs+ft1h2vcpkyU2yegA4f95sOEbfl8mRJrSjNVrBpU6L3HK5bRSnCBHF
RR07fBlTyU8YttCDBvrDu4bc+KcRcXjueFewVWhqYMWBjwXwLUH/qnTeWZgAu8XTXBfWBa9yQ50F
SaMBeuuzdpi8ZiuMuM5F3oqvbW1Y6akn7w1q/5qThqiLcJI0B5VG97ZX/zL8tErjL/CnK8KKtfG8
LKdIrjxdp6dTrVof9AHFFIDL64Od3uQyMjNTEjR3Llbxqynk+LhzpAyps6qBa2EdKPlI3t4THlpN
BKm3es/fXJ9eWLxcE6oYRyTc3mjQwFyX23cO1txe2jz6hrtwU542+rjbKfjydALMTPIIRE0AJ/QG
7DeuFcvTPwSXH5pFaCnxKMyXovwdheJeboIZUFkhDzeMClTz0FyqDe7kB3LIa07+ULT3sp4DV+XC
oyJJ7tb0KL+BtqHruirk//0/K7Whx8irQMCzj557tlvqNGTBUzubFk6nj2vbX/kmRc3EeJh86E2N
2krWjx3kXckMUfg22a5T0TPclwGlfOBikCM0N9vMF9xkc3gy07ni2ZPqOJ/8AFJ/WykVEEIpCl3p
nJZrZRwl0gdh6UJkqRCg4+eCPUFz7fTdAPBQsNkX5Frvvxg2RZ7MJ9WbN4179porNxGCKAO3F9tC
F6s22/YYVzkCNBnyZtFC0AXXrfKK96AvLIECBG1ScE4ZLb8wLbIlgb1nKyJs7ZxWD8dRnAMMM4LI
5We+ocyzpsUNgxzvlcrl6ByPHMvty3gtIdXqD1mnkFc2DeVafH3ANxVdVQ7FMdGaqPFf6QSxys7Q
ToiSDo9n0HYdSadQgufcZOskFjVBxud66pqgI7RKUmAVFtt6+uepjvi169lYB+Hd29n6Rh8+X0jL
lNr9keNrlu0w9kT8AC71eGdqyDuIeiHZZs1VygmFOI7BagS9m+D9LfP9LleUA9rUFcpemnpZyixB
EQXqvcoV5tziBz0QROlh4EfY8o8LgCAQcZtAYVRekrOw3L14/GY5I1ebOIoVA2ZAf90OO0H+gz4l
BxSqyfSFo/4NzdjsafYtvGOyAhXyzQj4dWRhYGrjRDgmCn3s44+2P4YP6cWwkBS/2csb3nhB/ueU
Y9r1GDNPjrLOoXBU1PdJYglVx7bEbSzhGk7PHqJS1ReiFAWN4RZo39pQaMxFYziDuowJ80AoNuFT
GvEKt2/06hNjVonCARqXvATaGdOcwwVH/LxXi1DesKVzH7DzFZ8bQ53sgCRLeXwaeUbj8AEXxXO5
SoI9atD9uM/f1ovA3u6yDY6gP42Ys3z+tpojHdKJVI06WGL3jVHifnJJyPS5TobQn5AFY9FVa+R0
VO4WrhIQaIsZEE1wIFpDvgc8dpg2xOoEhOSb35AKbtXA9XNdg4+WljQdGo3NKXJSW/ITLL9kvYgO
GVJHricIqKLd+qMR+QWfy086l9CgmdAWp7e4UoK70VZOSK3ZlnFfUPcOXW7PvlG49bsllWd3DgpB
LzAv5vIKiv2gqvtPm20mChYIIxaR8levwRZb5nNfFhIsYWiRWqJxGGQHUoxH5Luiuabi9L96+9JE
w8ylVUwMTLYn5SMJ5HKrhy7aACwa/CcUIOFt4ivbhKGR8/IqSciZP3PchGl7FEFmY/DRvpDEH4Ul
SXmS+BtE5lhtpVsCTrB2/TWQLxxlu13BOxevbK2rMG1QE7LET66CniUcL5jC5l35VR4e089zgsAG
kpUCfbbQCHncOpic8N8E8c2wplnhxxkyEg3X74YPN/xh0IBIMqmyLGzoKUTQ0VCzaqHhcHITPETn
sEMhwSfadQx+JvOd5rvUPr4gMEbPqCni3DFqcsQdlBJWTDiaK6HMfyIm+pZHiR2WHP+UxaN85xN3
blUB/4CWptpqKCd/8t7BvpUuvFJTNJJIC+oTMhtwNOWQOSZ+RRqLyhZOMpXng0qGo0hFbQYfWBMb
o4TqeZPKVypNM6Gx7LcFxS3B8y2SfLelwpWaaf8KexCvJLh4fBc0zFjpFZ1xaSH0vCkA6yK2vmzw
OzCo7klgRK0Oh1EU/T78XpxhqkHH3emtfdJZz3GGe3Q9N71x0TNyNd9q3sNZFIhiUwG+6BEX313i
rvRtkiatnhCulyU8dcKpTR0M8NP3RG0W+U8heMOSaDE67+m202w+HtwS+wT4K0iPNrh+f62JE2Hm
lyPDnEPmfGiB8UiLAeD5yjJI0Akcxst725Jie1O1zDEnTylQ5cskH6ejdU6BRDeopB7Jd1oN+4N4
tVALpr8WregZpcuLDOJ1n7WKqMpjShrw6QvUDcgYGrSaZAf9IZGW9yzK1vwp2k6ZMnWf3phujy/U
VxYg1RRSDxQPmCMAQRR86v8A5bIQtkOAgt8QuYGrh7KtKF0tB1AlUQx6hdqkBLQl55VpW7w9uLhU
rIsSExxHoO8emoSWHsDjSkvxvcoT6Nx4ZV2YIuvU8QQm9jTdKdAgE+F0ic/+wC9xYREDuPHTWPk1
6V5qiaDRq+f1wuLWTuCThhAX5iEFUj2Ue0Xdv1ZY3QJ/mxF0MfcF88s4qAe2gTMfSxBtkGt9zaUi
Ur6KrPdj7jLVOvveNZteYoNhdxBYoqvSO/EEtMV0eUaQ8leNYxKqKAkj5GtvDNO1Ccxp4UyhJSMo
6vxqTi/25XrcXDq4fljpwvsGACioFD8WmNEmnoNHVOW8fms1778608HnYZf0ljrJzCAfiOy7kMP0
utcW8YJvlEWSd5JY9T36W/Y1qFL7k9JyzgStz4c1UdEKj4W5GUIfaCqVOk6wPcDPMjKSGbvH4Cmq
T3sKBofmNM+n0sWWBxkimZ8MfYDg5Tyedctk2pSl4LudBgTBu8WYeUELr8c08k0uNrjTHBbmgLjN
CdlxgTatNTk32glehkPWWum52uWFRAmkaNdmYRbM/efhS3T10tDnx/qux1SDNTaqYTalGGiXNmdH
a9fvra45M66Sd77EQaXu7tXR7Tpgi3inyFNoq6miz3ni6Dnsm8+IrwryqFiYKJyfsPbk7bkI46cx
XN8aD5gTFTBmrvdy80mOqe5aWTmNwiGP5rfWOUusXof7WcaiR/uwAqWEanNpzkVKrI1V05zPGM3E
9xuQihEBhda2Gp6MSGih13iXfmjLOLlQIyqUEJ9Sns07FncQOTLyKIohvLMilvRnbqq3QJMJ0QZ5
inGBtO1kjm1t3Kw6RtkZCtEFJA0G27cguciXT5u1hLS2zvFjpbKLhnyYbEjDjLAkNq8vuO3iQYtv
gZGiTTz+T+a90xdGYDwtczpgtf5u/yBse0yTHbsNAALW6xuCyjTik4ytNmrBG1W8/xX8wwZ39hYM
1rvXJRUVlfpBtoxx9fz9Pi9eLzjnulXaIX+X8sXCfiy8nM1VKnwGEBjoMNV2ne4g0AFBXB67PtoT
oSWSzj9oy5DAsPdEspapM5qRVJSYo+HUb36WrJYwkiKdebHwF8mELCx4j506lHR856Wbn7t8sa4Q
EFjavj2bqIo8Qhv/0FWOklAFasAt33kGQ1P9tjOgsnV7ts/FdI4iWH7xoQUXipv4TALPcQdrD1W1
jh1ZKUZnQEXxZo9EniJEpXYsGdL7LT82m6QmPZ82puVDkbGI/UOnpw6WoNS644RUlSQNlPkeFWIA
6+Dz8SWzQM23eRB/Zz75P4uzcvf0pur0I0UK5qPZ+13wXbRYaT7f29c/VyNN/P7gkhZjRGzXF1C7
8MZmL9CeDMGTyLKPYx6tsz4Roj2eKNYPQ32F10Ll/2Tpu5N3UaBGR/VBTcTeCH9jvPOwPUj66clO
No+ZFf5X7q8NN5TD9FThneqw4VUSqz0RL9M+y7vu7a7uzeHvRb8gaGbIPj0/uz+fPxfPH+sJxVEk
Wb+bRmVEADJ+fL7rnlEnrUWJ+8I8XclfjD2/HQVrkFpZpFk2Fyeh+GYGpwDnUGyHxQ3JBrUJsKtR
YnCPqSS3k1XyKiS/NhEOdkFH7xQ36P0PlpxxwfIoGB/gzfjBXNwInfe13mtYRT4SHQqTRJx0DP/x
mcibCIYwkx+6pY/Rrc7iHeGhsKv1p76r2ByoI/vfNWHLoFRoPTdZLRqkEp4D/EHN+lBtQvSGIMJD
aq7RkNpKD+MZ0jz4KHtKSx7EiA7JIf7Vf4pB1IF/oY+Nw0RPiDp/McjHWrIiSMUX0S+08/T7WWNa
gTHMb9g2vH+wpk6r0X4LUg6K9+eabJffArS0OXTQoqdlwWSHOAwU+w7LpAOsOVh4Ne8NcC8RVMq2
pxSNcEd8RULsIC1IhFS+ppKkEgn3D7w/askDNRInLg4TIO7O/kEj/pUVXrZtimckJs+51EVnMvCl
KcYVMgf690Ek0//g7HjaxSnX6zZTx25RjKEkCm/P6XBMhgg+rdWpzu3dJl5dRKCg3he+U2hn62Xf
xnopu18hhta93VLAPXmOYVDE9Ls41jQg7d5N+2+2sjIyJ6YF85PB/pgwpIv2FaTDlmI0AgHmBdMB
K1qpsfUfAwko+SjgLsbVLX4ohA63ahNQLdtSy+19yOp+fLRXqrxb4qLIu5AyHnBNqEZefAFhZCeJ
Km5uzl7uxCaFZmz+ofddS2Myy/nVuQN52vQdS2I8CJUGCRfxd9/JonrMS1fAEzZ4qIcKfz82vrWU
viRNDVoGFsqjDoHvQfGklPjz5iWi4zk2rNDE33iGo9CZi4u/Pma4bG6KpZLysZ4ndujEgRhAvuFG
nRbiRXJanQtfL2D4bCxJpqMqERxj71sPnG2ddaEbXiQWxl8VJq56plg6b1FYYKwKV/OQM1MCj4qE
Y4/SjTf7OQjp8GGCawa1Gd1SOI4HW4O2RYVR1PLs8LuyjRjVQ+/fp0/qfw4Wpcd3+K+mmnh6iLY0
y+n02fcE8v32rUpqk8v0rFQRvJRbD93hwtXIPxeh6y7EupRRfPA6bg4qGPvJ7tO3acKburH9lgIG
VR/J0wi9PTQEqHgf8jJWFAc6Ed0R5DimAZvBG6FN3UckJcf3EoL0lHZhw0aniXh6fgfIlplXXIlm
f7Cbjdcc+jPjFd/dPj/C4KeVGhf7T4mkpFVLZYri+6+LBdCS2Lm7BhLfXmF8TclQquOiwCEzOd/l
fOR129vKHL4c+paNWyXxr29KefF6JJVvfqPVGErPYBY3a77e28BckGBBdNCxbGpyLj2kbFFhName
Z6zwCX1XBkQsfMvumzrRaL6dSeTjZ3lbiYXoSCYbHVO4f/mQHgTJBWkiioA/IxNLXLuvFqkGwMr3
QDx+yUqnEJm+tesgAu+QOBqX8qHDKcL3SUE1Dc2QqRABX0bLA6VWST7s7VzfrfDgxabk7d/wvCLS
Wj9qiSzkmnyJLWXpVDPZh1CEzqVW/f5mmRw5Af0n0RrN5iiU5J8MYEpvk0ellz843+M8DA6/g7n2
lGwx16t/spC7TW7S7IsqgzfC0tO0YmNU1+gbQ6/QS8FuyiU6+q3VdI/f8jm9tXwqIJA4Pg57XI05
9f921nrAdEOr+uPikn2pccw1ICBaudqFwnQbkXpBqvguvkSNFZHaLfNW0Hfw8A9c4UOWS8fvIy05
9eD0MERfhK8tYM+MNBxgWpeaWrPx08xoa/EbuoIYsMmckjcbr5FoV7jS+L6ra61789egrbFy028H
hseZIkyDIe16cTEbEPjH0sDQtCd9FYYYcHaoGaHoAdkLYKt9cVzC7miXNdLSjO8EHJRjqnsDflVT
z9aE+5M/yeCT8d4OKpDK1Lfa+u5SvlICaIeC7tW1jclmNsehNxUmOM95By3gWoheg0eFEkyqqADv
o/QSnNMPETtewBx4+FThXN/AxOpVbtY5KbhqWiUfCEfQ/IVk2TtNyfk58iKhSIceePz3rK3d0m96
SmH5f+79Ijcl/pyOI8tNNSPqOlD5GxUcv0+A5WPRAWZbpADacmFk0W82Wih8y/GQSVetNEaS6+Bq
znBfsoMZ5y4VumM/xJY0of+A2ciysaNYOKI/F+Vxww7vd0706GD1JVB2H+gtOMjcuwK13QvwVkXP
rNPIUI9lq0MYRoMK4fclwytDptdnoM0nEStFvfT6aTVmAGvU5nVV9v7Q/5bVQbSOhQAIrwA4F3Ji
qZVBEq+s7V7Fd3bxd58SMgynkrJ2z/iq0zTwvo95wyvUZCcpEQ5S4umszraGmUGQuVoknCvL7Max
RLSmzlRQMo8wk3SlBLTw7waxuJfAArZHKF/Q5eP88sdpc2hgjUIKRyOHMT6GmfneuqkPmI8L3egd
PHbbLC6/F7tWMdh/AShf24F+kncq6MYD6W+KUddFb0aWOfeqFg7UmSmo0hX4NGpDoaUvOuJjAVXv
ZW/zeRi+UZeFw86TNCjR9xzFZkyTDn25tZx2VHDkqq0hDW6rY79tp82teBa6z5j+cge12yFWVXvo
ebqhJM+L6Ar+4Ne7oDh//Ak8A9Huv06JK40y7VeVGNlS0PfisBlt23U7IvjQmxKh9g8LpowaxEMG
E55tQkBeFv/e3mOxFq0HpV7y2r7dzmPrJsr/ut+AdX04jnWFD4iyTM+xbSDcbrfaDYSMUq5DZkc9
7UgYHveYIrLFJEcnkARlNLIKbh1DAzxor7WuSl6R0jOQJ+L9IZiLgHED+M+AnaesPItg1XiKkdH4
VsKJZCb21UXkG4GD9VDHP1405bcnaGdRfY6VZEf4fd3xkbRPKX2Jaxc4flRP7sbrSQSCV7BmtVyn
Ylqc2RXkrflQ0mYzjbkKsUGwh4plAOgADHCV5QfjLhhQ3IygGE9UVRb4mJ7qrZ8JbHNo7jm124Dz
JZXnPLUPAhyuYBOFMVaMhQhMtTWPIARXWTnDDLUSYeJDhF33D5IhGG4YcMssGxXY96z7FaKGbDxg
V6LehlYAA3bUAtktbrgdbFnOSfsR5dKT3rN31IL9jYyYKDTv7Cc0LQS0iBqkEb2pa6QXnO09zHpD
8iLPSuA/qW33xYKmJjhLYd9/eAQFZg0r6H1ieJQ1BvbiA0aPF8fjbV3fRnuczNxffcSGUTSqoQ9M
TsxYSUcNaL/tRT6dzxv9sI8UEmpNo2OsQuYAjpG2Z9LXBolMqtZB1ZT5MHbJX9C2vpu37vf4MMp+
52wLo3pgqKR9GeH7bP+59LQJ33tHKsFuMOUHL8DwT4kzyAXWIPlewE4q4McQCa2GAMNFlWFEhZDO
gcc4Brwa/6+JCm+8lCIKitF7KcN82RSjtNGNgrJ0ARq8sd8j9HWiEfJc8z/gzZdnqHLw+HlFc9Io
N/D0VF3/D0myvqaRSUW4R3YRB0WXyaZfbGzwSz+64uC1fsNRqtLhQ8bDDACX5JWbS8YTaQGKDAPf
EjuLcuYP5tSoZY5JpL2qBcDJcKWZuh+mBXz5fnRG575hHWFbwYojEu4VGLwLwoJERA+EsMhgZeK+
GmJR3/ikGIAJn66kRdqavqNzXkVKiK14um/741t9FqXiMQngkksnfATEIt2lwADS+M819exrS0vy
3gUAVRhsHChn7U8hPMgZ/zF6icRVLwyqmSkqP6iw8s0BHAYXNK0/z4SAf90WSyjGs4m54ENAsf1p
eCyCwQrAvyDBqaoojkxet2K+OqdjZNzFR13s0xctY9nQQSUjTJ5vnE7CJTNrmGiw5Is2l9Pt/z6l
aOSSPTeIwZxB9+pUZMAQ8onweiPplsZE3ePT3aL364a8FD+xsLS6vCL0HKuJyr2Ja1Y196YfRvt9
MhbvdH4rMatum5PEVSfKK16GeWEauh6UThuiMgcpFlihD91Z+As/D8o7x39R4hFjBSm5+9B+bXCP
VzeTZXhzcqAKLKrT0bmvu8Ud2Fj2I7uGRDcEFRCw1BuP2rI86fbaE5ZGG0/K1KouTPjA+ohIXzYW
ZWBhV/yVJY6uCIolbMce3YW4LHvD/Xn6TXwbGkvBMMZq5jquLe3UBw/6elvpeEfD5O4tFkv6rXZv
CIuPSVD2bEjHR/VtcJ8OaRAWTGfGh9ssglvi/dltpN5/Cbj5alrleTGOoknCaihqTlKzRq03oog2
ARXh6J7Ml2WbRDHDKNk3YbYf8s0ByvEC9sZF45HEQBwIORQ0MQOV2O+A2ZiiiNQkmkOKqbNwf1UX
TmlAay2ipBlDKk1HctQ27Tf69APsJCyEQ1QGZgmJ4h2tLu0QPF//+DWwBIhDF9dzpx012AR7aRY7
LO5thvXm/d6MLH2vIaDR/Xb0BF0SxDqnHowy76oUAiYlQ0d1T+hASpBALoqdBfM/nhxUr3hAj7MT
2efwu5PzEjXWo3AU3h80dVsURh/hJqD6E+tmzS+XhjiLNm6cHNCJhzo8sNSKWZBHBnMqfVn/8dlm
8p0Hk6Aadr6HRqHP1LvUqKiXJH/12f8qk80MDSZbJzn1TP6tMzv+cM97Jd4dXnuahV0z1svZ3WFc
zVH4aHqFUrS+y21TSTzoV/8MKJuQuIAcLkabzKDcM7+qJBVK4asblIwyfcME3DUBLXpXSzoZ58u6
ZJRiE4250Jf8LjnmC0g0zx4CHcowbZ8yoMwhH3Scv/MszRGQKJ99oaVLx+fnoQAEd7E4mJfmSAsg
siUib9oO2Pm2shD35bx74Si6soBhGE2jd7F5EpKglee0XFesbHkHlJgua/lzd2umGOSOO55Lyxq1
5ISlCv9BcL/hlv7CM2sIQPH1KYbtC3OqGmT+1Irdl/hvOFuslVQDxTNKTMYgHwpfX49mIhYU5FPe
EDhz9rt3TlxBTTGFUxa0gGCpPMaacHpDL2fwQB8Dm3Wr4Ta0UClPQgh5A+RVWoIuXbDV7lwaszDB
5vgD3k5MnUfT3xI4aBWT26xRr9TNiThPjFuRyuYoun4Fu9+TDmwQ/t8jdTT9Z5i8WqXU+YYEIuTp
iCFVv+9yRsbaH1ehu8ZmAVQzr/dy3MRAaIM7YFDgqpyJMZ3Brh18RPCNNMVXyLcqDGKUAHizfK2u
XPzZvyPui9/iF8cYWc+MhU7qVSV9Bj1XpiJAGD4En55rcyMXD9vPzPJcYDmC8E2A/61ZmJG7bpN7
tpFqmRxsgt7Zbb4rvMCHOKGLPxLhGIV8Wm6j2+UGhnI/85YmOJXSCgRpdPm/szmly+9HW6AOA+2O
GzDStJBoKiq2uz1qmNHt5+KryojRwh4xrmwsy2MzDaAajccD3HA/U7qM1wetyYJE/w/hSfuXh+so
R6FS109px+xO7+JP0sYdnzZQf9luJOiaUtuMeejh7333RTh4oOwI5+Udd0uJjMigup40JGuN7H8Y
dtOxwi6B76otHmrmmMUuNTHP0FJ53ibD3c7L4CeWeIiyuz8Xa+nID3UFwcBHIggSR91vqEo4CgSB
oTFj9yNdMvBJVCTEr8g6l6Wu1gOOrv0F/R90XkJOPxrl2X/Q5K/9QynDe2+YGBJxx9WyQEw/Zxsa
ykjZtojfTZmfkvaiKIYjU8sV+DAd+nMfa1bRHN6S/BpIAxhiVgUF7G6x1aC0kb4hELB/Lgpd1vpF
wQEEaFifupigB3hQmBrNYd9cDgaO4PRTWJAIJTU5wCSYD4W+zhWzI4bb08iHWx29MbGnZAJL8hVL
YehXEjleWuIYOfA+YA/obrLZDia5JkMUYCucT1OxZfcxyvno8HxLzbR3JZrASKWY7xnxxo8e8bmw
xXaTEhkSknrUvHKBTncBaVSe2j9mM3v2q6Ql6oR3IA7e62QVQxJB8gWrsbHzIkFJ1qsuVvOLZL7T
zl/aXMgWTA9lYdm8xACzSPzShUpZZd0/C3IR/Bn1fy5ozGkrb4CfypcgMGL2H76ffNmacbFg3jDo
SAjGvcGvzTaqwokHDOnf0Xi2XQBTIjYrfn+q+8VhmW6k6KFFyPR2FlRK0/MsIs107oeWYXMsOfAQ
kCNMvIsC3NDHlLAGPp7HXlfFa9xo5yN8VAqEwuzPiKDzYMQuNK0Dwmczie2KioendhMeTKR6XaWY
eJBiIKcJpmaZa/T9qwyzyMJ0YsXPj3MD/4B49qNtv6icHkr/JVzpwsjzpqJMBp3jH8dxIbeb+FCl
BwSKhQSsxJO2xLkZbttB7CEaB001vER/00ZgLSGIPEoDHutlrHU1/bBfmW56TUJ6BnrGsLRUDa3c
di66vbBi0MLE1n7oav3/bsBbvhmNVq833Ir0XvBoI9fGSv4EDPynQMbWMSEVz5NTPQIuQem8DQoM
wMyJlzfw4jhQW8z2InKoqmIiwLiCPghzd7EnVsA5fHRxAvBMoWrBcr0JHggnjnJr0R3lBw2DK6b6
cnaQk00P6FUnmEpmyddA12UFa3+AWhi7WEuN5Xu7s/baZK2Om+Y9XFfk8jxQHBxtrUMjihm/f7FV
og2QYS4dzzYeAzuiAQZoUbYNr7BBNECgYSeEwXdpP20HmXdrknBrU6X1ELVTMjgHviB9HdgO2NgB
6QZCpCXbfSVfVfKi9hjk3pm6lNanXWrsWBL9qqaWryLgyFTNDJ0xAgVGhHi4QL8hWgE058XsRqoX
zBDfbIrlIO4ujRQr160K6S2LGz3g4E5MUbzU3dt8PwKiRysY+AlcBR/pI3HobFXe7ZI/oAqfvSCP
qm82d9pbwAnOo9fmCz1/EhNO0UNea5lQ1XPP0QqjiSeVzbga6PIAHIqw5JosCvpakkE1UGmJz7ee
IAHnYNoSpq16fc8PmcQmxEtYbNK2oJZdQxpWt9RS1tfP+W6A+JB4C4oawGxKDeijrkPgeLo5W8+t
4XJnBCHUvJHB91lKUaj80U/kfJvebCm/sS+6TMv2i8I1qcKxCODmjk6JSWVk70NN7NyJUiFlEiyt
cozCZAru1KjqwM8IjkZXP4O1VFoHBMyFRpAOCGndYQTHV4fh6DNJ5lrBCvFh/HUKVNLPx0pzU64s
TprhEjRBp1gG4Fi777XGewC1KbelFwWXZDtTuV1bYVqRFVSxJ6wvXqEeNQ28vF3w3xCmVZ412eSu
KY+nnJUC4yuov/Z7uNyVDM4KUXg3iR+ud1w1vE7x9kVzk7pp1PHkW2AVXZbBYFqGlAD5tiX38fV4
keWXsEQaw4llHgdnUXiGp9kKjmCYMRdj/Bu+Lc+ee3NL1ooqWshRiB1trzbRqTfwE4MuT+j/2Q1O
2mJRxhrtBUGmBIcYIKuNSogiEiZWvRcMM8nr6upvk/iODeAxvZDnj1CscuB6b1xh/MLw+BGBdu0O
iQqOhM/AjzL4m6v8oXae3rVbswLmoVNfmt3nCDuHE6O9CWPzN0vOBESyfcKe2ra+oxNtwcoEKc51
HdniWgTVULj/Mv4+UYsQpBA9SwJV9Wrl3agXLS6uy1i8unWFUKC8hE+G70afULf6PmuLrGIc2Lhy
QPXWpMUXEEjN58wBZEp5HnjkohIvfRXyytw4Lb9UTM2XnpTkaxqlnQETrEWf8x3CWJfQG325+7z4
epX0SsMP8hqaURRh82rSDO3MrNoHh4yceIa6v895nV2fpbLIx3Kl+l6Hy9gUHad+2yP/DGZ37hzM
UX3Pt+j1IVcvRcI7Ove67xFkMnYqoc8/z7yGQfeT/VyOOSNQPWV6zdC8yJvMvaifzy32jIDE3nwg
RwFYIkfczF99DeKgetBBmmdy9bMcPeAzfVGmDhk1miynTnE2jzCQvKyQaXl93OhSgnv1nL+F2wA0
/EUWdI9HQjDIyzTok+jFc275uebyGlzoEWmnyVJY/iWq3+v2tVpCbkQF0ZVIJBN+sabNtHzrsaxC
j/6LqwP+xgFEy0dW0L2YUkx7jX5edTT+Mvo9VjiYy9JfuwNZsn+uQjmTXrujpITj7Mlgvcioq8N4
SH7qVgUQfGE4LMA1IZdHNYkOp4hSXCc0j+YCQ3KBPA6yPFckUDdHMnwBY6FWiKE644tJ2DZGiRG3
Xe9q9tPVeCDxQP+mnp2zOSyn1xNHPfAzLgEGsAIURhqnwvvLxLf5gq7jkhvqWn1elBYpek1WF22Z
UPYO+Wc9tiOiylf7p1PM5Pq//RJQb0s4rxneqmvE7fsvRfyzo7tIgvf0VjCwdUaLIFIK2ZQl07Ip
JLcyySOns06gl5LnX/SR38ZHRyZ2hoVYLSfqsdGA2LUOlhTVzOBRLqnVAbGYqIn6Tv59MZW4jykX
sQXBZNXeIxYJbJS2RjfJaaiqV9C3FgQvEzfZ9/2h48KnfPPDlgCtFXUGBWgHsiWq4tmJd35YZwxi
Kje/JiiPY/DSc6JXt+QzUQhxQYHLOC+hNODjgrejInDNMdEkJR/xRejDRFZVJxi+6ZkCcWXLYjWQ
RzxGnNCQY8edHPGztam2qYL7InqO4ce35hjID46REH5qiCopLhgaxbKKJ7HT9KNmiM1QLTnYdGb+
Dvep8MM+JcmfC7vcZtkFsWtvJKuMrSGcstytVg3kKKoUc7PVNGEtTwactzivEu61qeXGHTJtD0zz
+Unf/+gydsjQbUbrSc8wWhxakUZLxK8xSin+gpZYe+f+eicEwGJ6VcIHzessTx3dmuq5HH6lmrOp
gQBWoebfuYXVSQKDd4Y/YmKKz38AxSzhpHGAvk5YUnPhfK/D8SsHZo60DSy5QmS0B6Vbqzj/yCms
w1ujjW0iewKdGMMkOK1uUpnPzcpUzIRBdwJxS5W9bTFrc6vmOCwo3aa4SUt+SWD67MADd8j0gcSv
BN6PdVepVIl+ixGZgTsBaSvNW+UlPfZ1EmmuTARaJdHQBelDSEmy2wMZgaZdtqjZrsVTP+J8pe8/
3L2rCeWdJNgKQzFeni7kvy4Yq1y/Z97JkHZOYxXFlNm5gBx7jG0JNeHDcRGy3e0A3NkCW71fUG5O
5bJdoU204hLm3Q59BWtih9UPa5tMiu32BCzEzcBWvD04aY9eBDWULazELvWQmYVMb6m3bOVOCknp
bJyTj8Pi16FFUus4njMILnPiPbQc/n4QArHJqSOpGvdgp2ywYNDlX4XiUl59E/MqkJuMZ35tYa7j
ZZasl5znxrImnK92Um1mPXMy8jB4EZhwjTW3V/MF91A+zGCDkGsvn7sloBZbHQUq7gXT0HgG+xNK
vQmQorCs8CV27BfjYIEa/CPXLUiJpgxh7VmmrmKkCwN+gubU0jR6JTbpw4k4i9HfZkeC2sAw9myz
lJcCnYV3oLFXTbJ3nOoWrS9H/PAIKglwqxJbG5wDtedAAftsNXBTwWoPJlGqrWliXJlwW/VnYb8n
ageBHt/RtRNvzE0k8IJe0ncE8jUETb+GJnVNXaOwlNiiN246kakR4biGovs/aXkTBzqEXu63OO1/
0O3B3rZyq+NClHu9VaBD0BuDHIbxY1ycm2Uk+gWBLRvgnvCDMY76tPKyxezz1rJXz+yUVK67AjmH
1iAFM787tXYiFAxLpXUQqIF4mDsc/lPS1IDKDVXPVh2AAQrwrPqE/+7PcWpY6I5UF0KBS5qU+o5E
UIzPhbU7TctfZ3codraQ6Ofeklkb6fDNdkts6bCeSb6e2qiDnjznxQc7jymcUNVATQCQg+mcVOzg
4T32P3x8RW+z5pP3qwhmH8bSk0pO+lsDpIgPbT7SAmS+AxfBmzu6P6DgaAYDrCC3zBunODEvjvuD
zYEky8OdMklwa2Nu3JBaMy2SrynTM1agwD0jMW/1das3wsIMCadCokTPz7taWhlQhxq8kvPL3416
ixPeI6sR48lyFkrBRLn8OlFbmJWu1VFKsMKLLfzxaGleZr3wteok2YhY/PgeH9GztViMCRXUvBpW
UCS8VKbMfDc+PphEE2BTk+GXW/K72t82Hosb8329VpoyGtKYw/mKPz9wbsW7tkkky/44/QZJeWJ4
/0ceAj9jgDf8HPO0jALjspghH5/drkXMbNM3Jg9N/8UK2eEk84KNQsie1cys6stVFC+8BS4j6AOQ
+A9QvjksLq6kmQdC+xDlgg5aiSf8JDtUkECELlw+xhq0l9Lk0OTmM20SliIlRPS5ewpQ6o1G4Mno
OlfuF3bS0c1kAjr9xyGCXFERyhT24r3x24+n3Ru+AUkAvJ8LoxyyNaWbiuWLjIAJ3PTISouqwwl/
AAT+VZhradc04gmvnaDX7r9xl7POa13CS/owrqejjItfQKwBeTbZtvSiFw3NURbnrsaABWI4nn9/
Iee2MFU04NIPAU31QRN12Y4qZ/5uLkfJbu6hbDf32e4SpViRqFaKXGm7vOlDMtlOo1aFPFvE9Ddc
zKZne4Im5gWL6Ya4/+ElzStSGoDgn/g0/MJpirgblMaUFyQzt6ZDdN54n9cp1aRoh/UqBL+pYjDv
n2cRo5D0GXDxdEXKbK04mQU9T/4gTlT2KNYjW3yecTi+SkFek9ecvtzP/pSld8K7ByrGncDTTDKm
0eejbObiB1qDOY4dIK5ay1CMbt/oVgwaQIJ6AjUOGbtXnw9uVDBqZbnGjzT4sDiMh5pbom+gKpD2
jZEL9IkVZoZC4Xxl/AmiUBWld4f+Lr9yU03GQWeMn9fEFVPYwuSXop2ury56I3rbGEd8Z/d4QVm8
RjDB8DBhwhZ2VHTeXwty7qYjn2VhxjQDT4rxB6hu6AOE2VqfFoDlsDVmadPuYX24MpzgX68Ti85h
UnaOyQIMQ4lTi1cuPp56ZaVe1+H8b8wIkh+aGNYHnuJuyLShmwO63800UtbUx+PdtdKP1W+1TvV9
I57hONABuwL5huTZ7gOic+Adma+vXeU0khjBSUpeF12zYFmFmKChkG3wLS7Xu7HKNPV5JglaucEK
QZDxe7p+7fM5Cf2rgSogLBaUVRmiEN0oyjxmp0Lf9bMffK0YmNwID/xESzcuHIKmt0gTaL4ekrCd
Vyfolf/4/I1w0jNtFrbpl76Br0N2caP4XO+qhANC+9wd5b2oyeWSYqLTMCZ9QJ3sV2KmVgPDziaP
1OSoTfzfszH77xBZWP//Y8dKbLxyoGuuRsRPRwsfs4/7nQwvR13krthGxFyLCMDzJvaMA/F//gFp
PGTtFDUVSiEcYTa2t03+On59KczT1Pyc5k3tZSTP8/Orj6ZEJmzrV/h8Ri8/ioRgKOVT52NBveS2
VTMMPfJeuFDc4YtHWJgm/AvbVAt6m17to+lDbKvg21gZow7pPgT5uYanDbTtX6RGzBCfTeMQuAiG
zBpHK9qkYY67497CD5BUWItjmd0NoKb0F/OI0iNuTGHW3RudjGUW8uRO9oynOs6Ahr9BiChofDWO
gQH+ttCVG1Kd4aXeZTMQxk2pLsaxucrG0IVWLh2CA6+qaVtwqfx/FpgW3AAS9UOL+86gxtSPG9M+
43mNpWm0OsxmYhaLyADKbDZCdVIBO7/YHFHubnirMZF2Jxxso65granTaZbgl2/PTbai9QPJuZdc
xVOOOLaLxfpZh3CRQOkXGdTxv+zZBKsU7Jg9PiCM6FQv/LYwkcI/QcPCfOZCspnI1Ob0hGWKMAtg
VvOqTZ75GtR2hPLRdvfMbhQj8wXr0IwjFU1/qlbmiIjnJgOygfH4c32gbkm80V1J0ehu8BwUrtae
FXyYECHVccEza2BBqkGU8zwXR7qb+waEHjzy2HQqYlHI1UDPVItnhFcab1SLYYPrWWJG5m3Qs+JR
nl7YYaqJhPS8VC+EAg/7bH2gKuphuDetLxXna//E/Oxcpx0T4+8a9o8MiQVwbT0usrBoIuVFQ+4D
EyiTAiHZ5G7vb2pqL6GZWFknE+kc2NsVu+koQj9zPdCKesxrs0D6qDJbE6B2tnUHzFT4u5PkO8i7
lszTIFWNz/QpSDqs2Xjfipmp7flHREoLiPxElOZd2UYs5KWvW5L0C3WIjFmDDKgK1b/nkbwnB2VD
mYO0//rf//+bV6JWK+5nmnN6DSVrJ4q8KFDVUptDKJsaWc2XfhTB7Gc4REmZZ5qozgkXhfNujDaS
HZi4kP2V3IwtYpmkShHWdiGu2+C+qkHU+jqfH3o0/YMPcFzLDuOzszSyJDKY8vuCQAdw6f0i//Sj
26Ru18jnNJQoVxsVcKi1uip1NwubCVwOpnwQ/evxRkWEaJYTTnrPz5UsJ2smecirjaNXJKHvlIq+
dnvJEVi24rgcEaiD0cQaj3dfOoXSJnuKakeEMicdbD1HrmVxBbP5dZ3kyhfZo6J9oX5ipB7news8
53l49WLvC4IHC/hZhGqV1dkz3xtlMcEAHz/KGat/i8Z272knAURpMTMO+7hwki5VFIJRPhdb/7ws
ZbBRapQHHE8taDIa1gso8zQqCSW9w4YnoR6KaIa5B5nNFhd958J4lsAxLXvxrnR+b0FUslb8nT/8
q26RQyLlErd381rG+FN1O2sqxUwfVHIpuehyWBjN3wnv2fn6l5iSore2hcWnl309kealLxJ02wT/
kXSEFYGTirduNksl7CIztyOTsd4dXgwAS48tZWHrvmrVpER0OUO0HoQcYD+nD/DMErOU+huXuyGf
XJK7kPs1vsAk/s0N4fqnrBIneIrnY5AWbnZC2sGsBO3PdPCqHiHafBAui/gCME4pdj+TKd137BMw
Eg2k/U7LWg0XjNe/ioc+XGIYiMC7r8V4b3zUNy7coIVb+n6xW82LE/UyxFSU7WQvlpNzuNPgZipl
8ZYIfrolLPFLIo7DrGoo6BMdKsKXxdqPiFgmf1PsmcP1/t9tNAXsrj5ApQX2iWChT0WELBFPALVQ
v3BYZC0XkQRPtJ3aVg5VGXs7DNLrXEgwz7nWHEICgUUJ9/fwEF64hROAedQHXz3vULl/S95c6KnV
o+ZbajuwGSmagTO3Gd2z7UFBhBhsDgm/7YcNk+G5/96CFsVTOevn6DdGKccXIUAdwNAJFpf5boHt
u4ZvtEvUNvMoDxj+RuxriKjbnm+9IpIc2hzZuxkSTfQXElWxGxM5n0q9XeqPGWiqo9XsmtFcXYBP
fzkwl/ekivE3AboCVjOlEmu1//77ZX8S52t6ZFv2oHJgFgkQAn4RA++vEHsatSqio6VOyYOU0T4m
eV/O4S1bwCW0iKURsuyBQP3RT26pcsHz31IGOWZfZd69Gk1bhrUHwIMTUV59vwt6Vwg0iTk5Cnz6
Tpxyi6uXcobwGnGPD272b15F9cB5MLBAz0uAhunWxqIXXFU32csvZ5Gc0hagQTVhA99ZCZsNsUV3
Nd4pZLxX9N7c+N6Jtqp8dSx0tEExm4eAdOmjX1eKpxu1TZrMEoQt7NlyWhKrgTwYesufJqzJHvCI
4wapx82rkOGfKgRRYblpDxp2aZHYeBJGpsaSlRMeCYFJCI3h/n4fywm7W1z0mf45QcaLFlKRa03f
FXw2EY72avUskOG9h9ckcKQP7lZ1FmCEt2U/76R4KSYVxm0Upa6XKEQtgKHG2ndpnRLWztA6sVTZ
ZrGrfk2sJwigMjWjzpNBRFl+RvvAbnU+d8M4yX7xZcUyjbBl5xT8FxE/kbLLNJ8SPB0C2CXRwDjx
S2iC/9Huwc6+zFVmJDLdc3PkUIo7uxRxXCKIxNxQGKQ6FNZonvpCuK5/RbMixP+aEwoTATLKm8W3
8daduuPZykg6HEcyKJ8ZDeLytdFOmznNuKzBiNhnLHy/n+qwRPLbXSqLC9azPWAaZpaYrZv66cCr
svxLoVNkuvVFHPxD3fO9coS8KpWTtR9K4TEUNduUbAl4f3AMCqcIYkIt9aQSu2Z7K9mF2Ib36GPH
18n3YvKnxtaFi2JVuXj/1tqqqCV4FlHmTeRwCAJUIKm12Ib90f7HTA/BR/F8ox4hThPV28ibb5nS
ouFdfEp6INnWHh7rP4CY/FGidizacdexO5qxwXkpfHuQaqQPzGDs2CgXGe73zuPxKsvEUXe7lFni
griGjZnu8ob0WpqUGcVs+93FgQSoBRFOjyFfHjpagWKYCwFbnmYtg7VyADZiRbop/hTeTBreWjWs
2acws0g/Y2xgWz05SylKb7IrkQ7FnDhgMNddDOtGTBXJmQR/1bOErci9HPrMOMWrYWg6yUySnN4t
FtT+AuNrxxqHUkwkrBt0xST3dR5RTWOE/fR3edM10Zv6pJxtjE4el2C1nFoktIWGFeZWNX7VpiIv
ydYcpgMjNgdfdf0ar6ruKE+z4DyG8ZSrKhLUId2+dk2mVlaGyeV7I7jzmZHo5f5ynO95iHEqqrWr
4nmN2XOrNJW4l1i1upzgcqRy1BiWelGPRXZFchLzZbBc6fSfj50kzuMCNbWd2TBmmqKse/lDPVVo
YGz2bQ8QXEso7zTPN3hx/q2c5cvRq978r/n/ucpLaT+RFR0uMMCf+2oEUeROcgmF8MafC/IoUxMh
pKkPF64BRBbvKJn//VyKsNl/XOZVPWKB7bVGA+ERGiD4InilSf2ar1KjdELnf5E3/7mOo6xqMlkt
o0Tlsxxpxr0puKJxM4MmeYGisy0JtRLv/3ir8+KGHy+BCe78uGc59Vm6tHMEUNEaNCJ+zxZIpkgQ
rea1CMG5IbdCZHceun4fjri4b0JX91XNAzhankXfNZWxBsUJ0noENAE/RjZUUSAGD5i0ZdUQzqKZ
nNE/WHy0+vaqCwYZCLa8S32c9OoTRcwejALtQHBenS3E5kWRhFz2O4DoxaXPCcd0OqpX4ra1ZPvB
F05BKyrDOMOzuWO5NkAGAK40j4m/et6Rr0LklebmEcawexrgsFTjDayxRjO9guldJ3K54hjh3HS9
fsNmzs/8KRklMF5Z5k1ZELsOXpE5FnBBtgGo3uJ9XCzNOMgX0IU2zL3yMguTxOT9pX+H51Vy4DK2
7DsA9UIyfGy5lOLLLGA3IOmawhXcvSBAWvN89NMwKJC3DLQUOrTtWOUCo4VHs1m2GIbVmW0xXLu6
zsamU526N2fe28+8oQsUPWqcnyP//Wnd0Xgs5VNOvLkoTp7yZMXZbeu7tFPJPCZ+P9Oavet25KdI
N9jaUkMLnh1/J4AXNQXs7cyOnZqgxzPY1QrWO9e1i3+Bmo2wmhMHV/AGLXpBCbqGJJDR/ToCMRxJ
GbTMtCEuN0YoAdyWaZQ2BFBLTogGjhwhp7aJFAiaO6GA0EmpsPem1tTn//4pPB8IkIh7SI/vq0mm
vd+ctBAGEYDWUJhuzneOBx51/VAM83VW8vXkpqeqv/09UXaTPl2uOR8no7TLiBP2+FUKMIOvrPeH
+4ZiAI3JKydG+t61wT9Umg1S3OvIHlUjzg9RDIgL8KxggnA+X6w1vBSpvxbCNg7Kl0Lw2bYzSJeB
2JBbBvRi7ibY2hipVzlHmPbcbaB7O1rJMxSvwklq0/dY+X3TEK/xBy2wrAZrl3p6jma4MbNoLd92
VeOJpuEWw7VSbQH3peVKXrITC7P4KzWTcGxDWYMfHdPgA+hFHzsdhptGX3A8n79gLMabbkumUhat
9absSsrG2jyOsPmZdqQZQNkRsEQzSat7oh/JZeFDQCwfKF04/+sOgwUqNoWf+0wPNqej5yGiQ4p8
/xSH4F3ZjLn3Vwu3onD4rNDxWu5oMxKw327+xbW/BYgb+mWk4skA/M2iOniT09z8+PuvOFh/1d5O
P0GfKeLfq5HnmrOBPBPn9WaxwWY1EH3NSftYgIm9T44mXqMokkcRf7Xu6YGzP6LqDSEENcviZV/o
o6fPRdS8CheJ7nwAUKOz3IxxDioXVwoWzZiquv3ZbNdKCSEMMc6pRkIcR+sU23Z7vAxy5Y7hN0A/
xnU+lTbnCOVUL9KFCXqhu2GK94MUyOeScile5L+zFQok/hAp1Q0Zlj85c2Tp+j7lCS3/MOBnqVf/
Fuac7jlHZWIU6DpBQwB6OcbUZj4QictJKQZwlZIQJ3+E+fUZmm95o/u7PtizJaJi/JM4KrRC8v5N
31FySEjXCEGvdk74p4AGYXIsyQUMdszimhBE9QvlTGRyu7L/F2bYNqEccVqX0lfM6BEm0iJfbcQ9
HGqqhWAr20tL36Esx2K9N0JXz0VIAg/dDDfMo6uqBVTfuC49dy2x0DtjITXTcVPiR40JSpSzWGdh
03koM9zy/tZbG6lBeAP2/NFa8zpBjErUJt7UuruaJADoRM9YH+FklmtbdDbxoQIW0UC+dPoKflqZ
UxTxYHNTpSL3Z8An0diM269398E1mVGDYgb7BAvYlUOrzi5IXM3mEWKcUVpgXH+YHNsEV/8D4UYz
9z6fs4cB6qDAkCz0m2G16fmPFB0x94W07oDSKA5OpEP6PEsvwNiGt78Pf40Tm0BtnOHSzrcJuNf3
fcdxbvelUzqxo6g5Z00ncz7lmOZebqyIsA8l9vFDFt5GDZEEHcS+KT9IDU34VOFaHOsOIRi6O5m7
XTX7TJGrmMxenlew0pPzarSjLLLFtKdCMNVg+GreBFTkbEp9G8gmKKtJ2IHZVHKwFc29ZL3dbli9
AtLsFy9p8juTbPoSgXsiDnJOPJGJk0h+3zB/7oQEqmqWt+ReT0epYttxdUiEbdEWVvlSu3W6kxcc
pBhMnEl90hxJcBlbi0IBvoqXGoOQJ9SCuFXIB3olnpg/bivLKLF9IGSwPD5Wg/RbkJndp1txEB1q
u8V02Ht1R88qPeM7CVJhUCLGHhLF+WpLAq+UVmNDmhtCJKvQzdfYQDXE/IL8h/uT11YvJkAvl3/l
TMd98fbY+Jiv00wcx3MjfeYJIvElGwLmW+xfwioZOwSfvRQhcJM1iMfoQOdEdjDlInFS92ZJ41G5
LyKHAapYDR7WzbF/Ab03xnZyNqhdOhbMvcrCEUGp3mPmejQSd5Jiy+ANUv2q3PmaMXofcW3eHmAr
KM6De25U4aMg41Een0cP83d0IRyh16MEpdcL9DacvGf+EuRvP4Xn/ACAahsmvpPAq5ghNd21tUG2
5FrwAbQdluSLNHm4nw3VUxRz79Yrp5BWl+LKiMD4GNmTi42MqUihTTiFsY4YgeY/QaBexDRt0O52
g4YP6aDBj8LH8+8ify83BJkxK/+Nz1H7td80d2tEPDnUe4rIyp8kYPiv6vumky03k0Ze4WQIzLju
aZ7nuJFwwOl7FYTKt8mRxwE60tVO8WILd0P5B7ZMsiFm67PNq1Jl8t2Ppy+p4Pa4ufsqqnet/Qc/
tCt0IDvAbBDgn4duMJpaKLpR1UUJBZvAoz+SFg/x9ZkgvrXdE3CTwZZq6aZN46Od8YbLIap9jfH2
xhJCYC6iC2ikmjhiGw1YeQPM+hHd9UlalhT+6cb66EKrlGQhMBl5ppiA5afJSyrh6cN5ocINgweH
f2Ozvkba6iEzHO3FOdOoQm6x+HgyZ0CMpBxsHVYn9F4m8mYcnMCkeneSZzSjkTQcdTBF2djksKno
+PNy+uRZIUG/Jlm/PFDoWOjcd7Clec1LXBbUChnNUSu3xXhdW4BMClWx6GjnrGO1pO9rjy6vssnZ
Cgdk8xv8OtFJFBe9gtnbSM638vTApW4v8J1wwxLy4HZPe+0+2Fv979OO/PvQ17dWjEwJdP0aABPq
UMvvDLLukR/TCKW9rWCspKeWADmrf8xCgBBkXgtDaK+vgmqCEE77Y74GijaXLOH2BBwgJRkFYpbh
ncKJ69PvhNTvNynSmYA9Nayr1JSLZq1SvIHg62jBO2KYCCr8MTuqsJNVpFbU7sr86cN4cuembEKf
VwxnvA19moKy5jg7cZuKOFj4UdqtAkvOOo7g+xbx32wa9ys8+L0R8CNIQDEQcB3ms38uJgI+LHJH
MSXQx0zPZglsytz+LDtf8z8PvXQ4NjaGxJmojakKdhEYbavfzAEnDIHP5pOO9K8agcGtXuJkc5Ey
N/jRMCpbTCN/0D9cWtFxQt3WMFPJQUgtZlY0yJuLQQEoPzMAHWTRCIHO7hpNVhJxBsCQbwjxCsiH
dWRq4tPk+g6v74QyKKf/Cch/TjlTCrEILfEhqM4iquTd62yej345mRSdDhHSWB6Rr+J0zBmC8iSt
DTvdgtAZO1orTtZoRLrhFbXyHa950k7drWIItwm/HP5URW8+48OhjRP9J2uQaEShYjNzWEuvrN9n
wu/NM3GWtW93cRnOaL613nCh7xzCrEFU+jLRdkY9bzfPh/N6NbQix6N4Nic8xsIzSWLFqDXXyq6I
8SCIqtgl8GKW4au0W+8UuTnsejPM0j6OfsMvrr0yJ08THj+eP03a7Vl0H7G7s04w9F0kEhOv0yEb
GiOSCZzyck+Nxi9O5SOcFB9XhnkLLSWZ0zgNNjbtoHs2QV1MQt+N5aQznwpLSi7ZJOtMPoLs2xoa
9oISIkkDJgK5TOckGSrrzWWiuD1koRyA02VrZ62MmBrZJ2zzoqggmkTgnh06lCw/d2G7kfbSWFGf
fGuw/CJs21GWUzDODDg/tmNIPqiIqsKZOhaQIW31gU6fVYOTJbOLYn0INNeMVOMS5GLmB08/lUNu
72MLH7UknuY2oOsADAkAUCRuPcbDkfSQi+DMWjNvYj67k7TI4etGGtZvT/yU5oIf/R6b/uiS5QsK
EGm7GJKMXTQ8FjbHK2LDW1QivcESHY/8BRmOkTJxg6NyM25G63IssgQTsZyDHtHzH2g9emgwRL0p
HSVY4j6TR0m4mM3aekdSiAAwz3jCNdCYRyL6sWEFPDsPnw1b4o4auhE2M2ybblUoQzfcdkToMrG4
iMmrQkIM3uy6+3Mh+ojEjXpJSwDJTs3f5iVSUtAcAFa/NntLSFWZ+pokVz5kHPV7+6nvHlzFsh4m
D1HurLD6kichXQ3S4HUJYmJ0loup2UVfwT+iG84wFUNqFJigPbxjCv32W2ZkD1ahGb+0sS8N9Lpa
rXzMioxhZCImQgx3O4fdA1btbHghzyw0IGuP/O0pENcSq81ILlVjCM6ZSL8zNaRffKrp35bJi/lU
hkkcQZcjGlmQ2lnGYaV/lANUtv0lhyOEEDF3zFk5BCKb29dkujQQGxhTngz6oetM5oSA8eGJYQLL
yW6q/okgJRROTooEwKhb1JzrnLIEquTHgCfxj4ahcnceNFRevOL521B6ea0vU9CVNwnKvwF0Kdd6
OFRWA3YkgrllRgv5VGdAjG77nYn61CVERSh1tFigWdy2Ln/mKKM9D+XvWtMT/oK0vZC/GuM3mLwf
gXM1J6RNlTRltR+QK4ky0tD7K16OYbtk8Ee1OQLB8u46gWhWZDkkfWEoXIHq4e0xrAfw0x3Wuuxc
UQEAfg/emRxiAmhPmmewVPFmKSH8dMECUO7K/WbnuarZA0HbRzsTVaMaCfwfB4n9zONdA6PdlhvT
nBpbaBI803m8ae2Zb8M9XIt2CGvG3D9uEFfSnsTmWMucN2mj05u2JH+lcZ2p6B9G3Ts9Q5oSSkz9
UCX9xStXbVj+TSVBQsSjABcwTlQO2fjq5h0pvN0V0t5KWwbI6fky8o5LymTcUwO1n4kaOp8Cu8TK
hzxIhZEfprV9msnfmYU/DwrLZnbc1DqZg2hZjlaikgoDGS8Lt2DQC5//xOOtNeRzIL+V/e5am7E1
wfNQ5xcEz7397Lm4OpGThUxUq38Q9B+XabWQkCJziL/Eg4wA9DYPHAjVQMPuqfUfnT+j0ANCxufq
0M2ixjZMQRc4LdZC7Q4zEydz1mOcFlc9dDJwyKNIVCT2mf+eFJuqjenhYql7h/6QNHhbD6nqsfN2
Xwn1wqtdSXJZ1Gauc1tY3zEevKE12hXsYGoUB4pzAfDDvLCu6w0u2L4/TTwlDlOvJyJ8iDcVvvRn
sV00yxxPCIsM2o/PbyDJ7FqnVDELLhX8VIGmJhu5CmrjCpRx/ZLTJK8M4dJEXsnIeAYPehjm9/Fd
6FLPz92XmzcflIEhn7BjwHVyIl+sjXya5CSXC8XnAFGyai71Omqj3+uZH/wejW77A/ZGmGCUEK6d
cIMbU19WQMw3BucGvS/wj//o4nKJQDhHwuushN15eFz1FsszncG7CtiW+oHtTRNTiNh7xZFVljkD
kIPA6IqlGukwDfZhByLNgrEJABfVklho0qWsPWwlwpmeYwo3fzWhSHyYDJTCpP4FTDgKHmEKrgln
3A31PPOVsZcHlyI/fxUBnI2qr+KM58B0nPKpXhKDMxpev/hEdyAAhHTatea+T/y8j7Ot203VqoQf
7ARqSsWsa1H4OqhkNa+/t9gGzyPLKgFlV0R+mA3/qsFiCw39NphEwTX5YhEbWGxs+F2AyLNsTvPN
l+PRRAzYFJ9hQLiwQEtO2X0g0k5vQeycHao8m7Ln/kmmFe1/FgfY93E4x7d1hTSZEyvBcHGmO9c0
pWFUaZGp8pBPZ9c3r4V2pU2RHoZjHEGQzw1aUS55xISkGZg1SLU7HgBC/KKJKBE00+ZxgjZv+ap2
1jxl7lhcs+/pcrka1UmjQP4HIubeR1wCHtoDEk3K69rQEa2QquCfcF2kZSQqFvFoEJDnF1AEwS9U
Atzj02bDmefADTaa+0jIdwgZYlqyKp3Y8YRutyQjiDDWkhNL2l+cNy+TNifNc+sSoNyTpGpqAYvq
iO0kOOOLt2Ixs7IrTnPXH0dN3SOP1bC2Qz9wtk9xW2ygWIX8giOYGtPDSZRd2rLH7m2Q0ufOw/pr
SevKf2D6FoVAlMdwWt0cRCnnpgZPjme0Kkckp0NevEGI8d2+lEIr3QI+vf7k7uThAZS00dPjHvg+
u3/dAhD+fyJK2WRWf4u/Qq181Nh0j03cnUJu16Cu9CfWEqhy3Fwmmw2SMwFt6f9KE7Lxapg5bspy
+8hCSqDLuW1u25YGK1LpVtJsQ1rz9+YnjYUq7JzTevN5/seTE26cE4PFafEdOF+BYfY34YU/eqv3
/kaTq24LxgP1KrPZ5m1c6PDuFH0+WHW1fRIO4M6Tulb/P8aQxHagDErbGrS9n6pkMVT6+Gt0KFJP
1Fh0efc+5FQL5/3yUsQFvMQQNwvs0YGTO2aGPuH92F6iYvMghJ9xWlkfnKcQgRIViA9ehwX2TJ3o
F9Rg+u783BiVZjBXCEAryE/bazkpyl3xVyY618PEvVgeJCHu5gQCiohpuOgNAnOfMl2oRJyL214Y
IRhODTj0PE1inMgsiqE9kxMthWybW+6w2E0d7jBbc1Ywq071NKIaYOLoVSiC4JTArMMfKbhZ9622
IjSlR3U/3YBKY4d9bJgwJTJdE0VYKt/gGNO121tfd3uY8Jyil+N6pILgbMVy14B1p+HsdG4t9c1r
bs7hTe6ToSmQaYj29DXSBZhpMUdDuQXrCiJuxxc7U+N/NG+qWHMzEkjPn7WtzudLcOopNYfU1BdS
8B01uNK2P2KX/EbMn6hrZrefBdkrjNd6Pn0sekrNWWYh+NHVHeg8IPpVaLeCn/44TLcj/v7lAsn1
uV+2yAx9Bulm1MWQ13HuX0rOKvqPit1VF1yHp1/dpIJa0msFNFhQVRNBL7xglHR3pZLNNUVSiUut
E9caCbtE0mGT9JlkWAZasyvnq+tk+bPTqS1Q8JfpRh0Dr/+WmiKhLXqyBDRlMkdjG5QbzL+6LJSA
J94ZQEpROn1wbxxLoHdEucthgYtebPH/Me+Q5J5W3mAKdfCL3ysUF8rbk7lqsWcjYiyCH0ScUSs6
hfamuMw7XZDlhWhqm0xRY8VSG3sR6aWeUYYyUbZgKquzwgiG4/uN7BtAuPIuiuHbVNoC1ISFBoRp
ZTyKGup+Mst9Fv7wba49b5zvTyJrP9KUBG+jBwgGjVMMDpZ/sxtRNvRlKbTZQYXzMOPIeHo8UGHq
MSYslKWmHeT0vVrLJlEiriNJtcitJUzQ2ae6Q7rrbarWxj9rTalGBnEcLUienpAE6ujO1gE+cxXM
U9bnhoNRJixHwePf4E4TV+23fKhDC9mqPH9Bc611q7qiKWgZgoW89HjkVXMk1lBolFWwzHzcoN//
DULBk42r7u8MdNwUl9Xx50Jhjqv/Mjr2c1hpCtBh18pDKXyal5fJzjQQ1px5e7VM3LLwWv1jMQeW
F/yatv+py/qyq0aMeSddhdvzsCeziR1q2ZzTbfCi1nSeHZhgEuAKDYag8vawmIl3+A1aiaxuC59p
v0Tw5oz+yIlh6BVLFBj+9xsWSMdY+wyAnOoNBsgrM9VRMVcL8jlrfe+1zl0LDFVilPJroxc04RwX
HLqeQtwT/wFh24/Pr2Pt8TwRqb+rFOlG/M/LvjkzIAGCh9eLgpEzHXRSRUIFQ+2ofuK/n6SJ5sV0
GYWdV68ICGh9WI28pP5Si12hl1BWeux7zg/LWrAnaQuHmckkvqZ1XEMb2C7bSn4d9/L/tOFumuqj
00mSvQZWu/3/D1XQb3aINyVbnYQUB0ZHUER8gvRSDNHDG4ox0UbvAk3JbvqAmfZpTNxF22h/bZuR
yevAKG3C9H5EUEN9c5dOb1Pk+kqMSvXKSoiFrFJWlJ5o6QmOrpO3/JiWxvFO6pss44Wx2Qfa0DCA
DwIVDuaZtOwY8xkhVfcZhy2weaMuR7v56AV2+8graf6KEeJQyMPcU7A6J7dGZeWKstX1evyimMoO
JZJ8ZSNihWHTdhPwSDqseEzYYRrXIbu5BhaQ4lRsqf7CfW9c2b0g/I66g0zJ3Sa+iQnOU9qDugc/
W2kEsXJ+5WaWNQ/CrbjOCcX46Oo5RPzypgL3TT+HY2H161/DQa/YRjfO+oThMQG5gjUccceLd+Cw
RgaqwC1HFVaE8xJTG050780YV++ra44jOUx74IWHFTpVdgxyqF7Z9GQFi+o/4GOBB8a2UGsviq8o
PMhln3qPd4NWkKL2mTwavA6h7yzRFtYZhCRLGiFQB9gWc8GwGGe+1m3bvx5Yosg6i5c3PzwlEFu+
Faw8ipsCBEsJEp7Uew5FNP2OGU82vF4Q8naXyywKTHZwUrL4me/zHOjchSd69sRyeC8TClMhb5fm
N9V+tQm/rkvYnKY0vXGI1MHLC1SpZcBckWnUiCK5yUbjGm9g9+ROrVyvtGy8npWeiG4qv1cmbPmp
bGD5DArtks5Q2y7RupbOxgy+iwh505NlPghgXfJMV+Z5haABz31Rif/RbXwe/nlaJ8IIKK0e6jmp
5XWTIMbtcqr7ceNux2FaKQR3WI4/+txO8oY34D1d8DkLr24If7mZNTmxKllMFoiFwQ9VRAc6MMxt
g8v4jNz5YmUhkYSHEPSpxfEUbBgIa9Nz1NEstwF2FiDteU30RNQnFFIDXFjkkwNUEwTRwfQdlTZI
TXb99unV0VNMvvad0715xAt2SyNKlNJeFVpSKf+YrNeMu3rK6BPMDWXH3L2rFyV4QUYDuPwTsI8l
++iEjfy5hL4JygS6zCxuJTD/UdwcEFIIwILxWhctz73zE7gHM2OcGTq48BNVy1fLXWnpC+467ADO
pjCj6+JlDak2tvDign+tDBb+4BGPJdEHvNKw8MSn60PLBdtuYvuQ+xo/tXU/8G7q1hc8GN3GXIVb
eGarfxUQl0YwBCkDB4IQSEUXVXrogUotYqZCVtYCVa2MuTe6lBkEc3YjhI9Hl+6UFTgewBcB6nLw
iJyQbNu2uGWmJdIvr9qG8K6CY1RGyhv+UT+FUYzJwmrCDutigqu63HlfE8e7LPizjMYFj0JVCcig
pdYT6dXO6AttQnvmJSH7tHDjTeW/G+QWrXycLCk4dCxV8cyuoPVLt4qxr8u+0BOd3+Ub/dklVbZY
JYhnm9nP48CBjp56ELX3V56f4dEs11K/c2zTjnHuAmga8BVLffeU4V6NqdEqLdaVNZryaAu1t49e
7676cJP9lqQJU0S6Egf7ALMhAu+zjxmHw5s+7ocuSi9tsCZwZwjHcOfNGcxRWW7+kVNjnhuVq9+R
1+xeBjKEJVrzcam4Rem3/U38473hQmHfnKWo/zBS4Vam4d9CUUWqgc5qkRReEXgPTdt2TmLD9y+Z
pYPaVqIVeeAVq8Ys8brrIIUzE5vPpW916AQkAntapzYU5oZ3IHNI/RpsUce+b/Uh118t5fQIDdzy
Udv8B6wHOHZAYj/UJZ8uoOm0x1cfZvv0MGFa5nzVjhKXNEMaJMaB5l5QueLDDt5qlxRsQSzeJI4/
1jpo8oyh+Ykkr9b6FhRY/6pukeQdkfAsOE0NFh0VVtHfDBOeXKd6F9DikhB5AUtUvlx8ZB/7o9MH
/qc8nxzuuNUmpzZACBLrdExGHEF10X/y+I0w50DvNwSg6enqN64OSc5NCOUDSNAfah1pFYroptfV
4OLWAMJJwTszCqsQmDjqexwhT7rKDUzuUZCuTO86cVNho9hQ+yZ+1M10Kjvuip8hsMT2pp6009sA
kpZrSctXQvfyDPliCanmLRR1T5OlOUgHeJLHxgtDQPTeNBeZW1NZwhYJ6fcoBtDKF+RfkPwTKNis
LcPptiOp5HwrNNoDyQNO3PMs0XYnQuUt6oEgA0iHmx52g7YoncjV6PDvUasO7DIiCBraCtTvGeqQ
Te4mnQQTlKT+l0/MigAjOK+KIuCkafPnLQub6vM2o7XpnS3JvTOTlBfK914heERDSCUy2LlMAq+9
6ua3dVrspQv7fjU3yE+kRxdn8GcnwpsQ7Bc/HskMB/2202A6DZTU3GGDD+zgn6RnaSGlNnXaiBPL
MeY07HaJgecARjMT+7wRL6jVSx0qp9mSFjJp12CWBDnxihlM+Um9sQRilZmJJpvhBz1DTdEgwetz
qzDwYeim/9AQJ8hTauLWDvGIZ1L4HP8w2V7XTgVPMIcL1XwNWFoT68thKGEoLPmhzFS9Z/+Alhvf
x4RrIdZUM7LvsEubduhevsR+hK2T07BPziWaNpfmWWTRp6xTxFLKaXxsahoRwPJEWxC+4bHP46En
hNDsQWNe8TAgVy/3H0q0jmPZ3kSt27LWJd911Y26bSRUbGzrVDo/TD7VGrUo2dSxArK89LVQfELT
x+FX/d58oLUqh3GjOD9WLNkKJU7BpFvwh3cbfECRIF1W+hURHZapTBlPoT2rVuQhnTaHuCcysWnU
xxIZr0TlzXsu79ajcIB6hto5ywaSYfTVGBwiPyLex4QDJKDP0LTBdcS91A/lRFP+YIMptwSQB/w7
gmTK7TXYwI7oiyguIRCxvCFPnpRoXYf4H7L2MKg2zo25S8sva1GcuJM5qLbWuWPHYSHXaOQQY3Um
dym9R3A2LNEhoPai4rrjtIn7Ri+UlOTQ17WSzRoZz1j4Ox18/wE7rYXgr/5NuQPcinmxSmMc1oa8
HPOuazopdhpz3lYMxPIakWqRBoLyDqHWkwf8gvO564PjTcrgt4a5CJQuldt+NagCeb5L9hMDn+Tb
9WOiUoNBjAYBdgGe5uLWTNzXdK80RWRAmxr6b/5Y+J2vDtKZtwqokYnssoFoQG4KG4qhp+vypF/P
PXvuJEixGYERJomow6Ke8RYIvcuv7S3mdn0tIU5POp9BFuWDnxraSI8TxrdUQAfWqs/lK9ovpVFD
Xl8GQBnxWdMzrQD35z2F12B2WQhVrDWf+NQvIgTDejHAO0M99NNhktxmyvHF0nCWqhjgtBFQz9RX
d465drfwK5FyPaKSuURIWIRQX8grOSbeE1lMGSbY7FNljy55rbCbQLVExnd5/jvCV5Ob8hxiMLUh
fsEIFdN5S+5yJJ+lzenvysnWqbQdlluej9a8oczoED0xfx6efBDM15qFknqV+cTHScbvHErlsgCR
zP7b1UUIYF2qt7rZ284ykZdbHIJciy9yee0emJbumFDTB2Br7RwW9GWwT5oKm8sMlGexVt5AAna3
Upj7wujk1g6Dd06R4bLyk/RUAdDxtVwuWzMF3IU6g8Vj8e6pyDzG0NHrnb8iIn7w3g9JAsCYrh9R
u56yeT5zd5jJMvRp6sdjhpVsaG6NIjtmn7v2ha+OGbTQ2UHuKl+KPe6uXCXdQ7lWg95F11EAXyq+
iAUO71ab1mUOtZ1LjXfa1W02Kiii0OxKKGP15rdBBq57Z2GhWCJbA7PRL6MgBSLlz6DkthKeEpmf
hTYXGUaQV2vzurN/ykK5i+DCJ41nGAUqJqU/aayASLp5EIzRmHw1PDBvDmzL/YE6/c9nHToPPHmN
R3j2QSdmUegVdnDsYu7qNhVG1Esq+UdH9TDPgXRI4Z3sW0eU8Yny2Cdk2J9v6GJcci7PkHDwQmsL
7Gre/a0eU3lhPaCo7LOB+wpbl5qPl2aJ2nKV+4PriZ0m0PGUiCdJTH4nMUtVK/FrRp7sqMFRCJ+P
wSRsu4qMp46nLSQO3AcFdtA+VTQVeKdnOz07X7FwOyLNpGAbn+//5bUCyJh9OUNOAHDbpcCX1CJc
7/ab8PFDPJHBrIhbT36u/upcAbVW+V+jct5M0Ut1ENQ82fHYG8SNhfSOBR2Dn8Bwd64z0X8rgBP5
GLbgx30wobxQX7LO4H7oOowAYgZS/chxa1so4jDfN8mEj8T6ZkLRmqEnlYxQDEAVFGVMOQoZRnfG
C8YWQG9lagU1Ueyd9xD3DSkEgB0lfMUPzd73YiXGrzq5ll5Dds9tYwDYJn8P72c7YkGv0Iukn8S5
8KQuGLXBuTtd2serwlG9zDF5QyLrh1R2r63FtsLaUmooIvOHrsKNR56HvaJrF0V0Z5eoKa7TkAt3
uMjNMXoSmf93OG0qBlbcqoWlmlHdMzQZDiMceESu0iC0DmWZfZrny1C02HVhg/Yt344qqsWAPXkN
jhsjOIxEGnWXlU3VxpZrGfKeEeZ3pJUODqWSRh15Z/CKZgohurv0nlSBReiLNTslgqQQZwcWPZaL
i/3FEkRtS/l5FoAktjFgVcJBlQm7CJ/8s2NqM5O1p4tYqBYtuK0xT0TQ/KIYCFvlYYYLmPeXtvba
75yWrxA8nzfYG6zcyus16X0cwfGoAIocFR+w3aXo42LZz/YMNkQsQt9clit5jLfBzIN8Iwmb6Mn6
Bza0WVJddooRbajHroAJuWlwvzFDD7Uy7fGX0e8S8ANCSs2UBE1oZM1tcAwEpJriTElPUQwQXvcA
lfblDIAER14+tYWUdUYC/oJPf6OV/b12yC0VU2cv32WjZeVa44wM0yxsi26RDBokerP9A/SIay2l
5GoeEwtoqt0vrsmTTbJ79prC9RC7wjFJmxC1iQZvh0gxAL0BvMyXwj8wlB1D6bN3d6aenPBIK0J9
R+HTJK6WFPiWHKh8EhUAhika6jBmV1HvsDmms/FvXGlrm6gNYA8dZiTzpYPJIeK6CfW2pGIjnVRa
luWyklHihlR4OuTyRTcC/5kcM5LzkyUijPV7tPxI7GqqqzXNhqHEo6ygPUQ/yX5wkh+JA3pf0O7+
c6DBFxzYuXQneiwPr/AzLLI9dBjsGPePFfetKOziivAqvKoK0vBreByaJ3r2lTMuZxo2RkfMjWUA
Mby2TZqFsDp80HVzgKQAIf32UJgzZUgo4WpbwXwbKZ+189FrzEQ84mILKvE0+SOEbyOdsyoBJYKl
d3Uz+ILAnzttLqMWI9U6Cq6eK0yME2FDdYbYG/gJ1T5BVi7ZVTPlsjnl2yismkFuEoXLqsjrjDUn
bge1CI1HSgfBmXVxUG3fXhXP4KS93IpV18FRqyzPtGVdzMkVHJatEUZEe7r1L+m68rSJwC1G4U1e
CXSf+s1RK1GyAc9NF4jpk8QXkprMGB6ksOrPy0npQ4oByIco9ebnBM5oZbGIlaKk7LwWH0t7xZTS
AlWQ19tWOfUzAhT+5Kq3z34qbs4dSr+jZ3wyiqZUVw942mKg83264bC1Yt+Vsm4t6qgb2RsCk+oj
Hd72ERYbxaj+KymSaZxuI4l5OJ35t8i+TAx9GVONSu/g2daISeD4PgfTOpFPtR97k0US6qhRowlJ
1HaM6+s2XTAyQpPDO/LEocJjaG6QtxQDuKDQeA2EaNWv9kq7dOAMMdaJ6LLTX14Ue+nzNpsXJdQz
P33i3a4eVNCAqUANmNmotqppTGIf0ALJv9Bh+IpwBazcyLbY6hnsfupbUFtt29lq0LMtA0hqqIhw
4DEAZpqfqtE5kmhCKOsXmVNgQZzo1wxbjEjfg/psefMDVuhQrfmAz9Ia+DUqUAbAWURarQKwV4Sj
WeG8F64Ezj8LB9XStMhm8/s67BZDVKxq28tZ06xyI/xN+PSKetzinqnwQiaP0l0/mHLzTZWaqIL1
fy2oJBGjbI3Im/VVlQm4g+bEHK8L6Zp1QP2MxutNx4s/RmZT6yu2AX03n33qmjuNxWvU5kmelrZp
fNkQIxBbqbtmE5br0u/AdgetDP6OXoV7sk6eR1rZ//3U0L1m9vO6+Eu3uRt2J/hwH2Umg9ZQ9SWN
B0ndVb4+b4Xgswh8k1dXPsBMW62KhA3k6YFb+TQt1umnmfBKRVPDdY9lI2Rn8/JmOKMGkc+T9zZG
JXnQf5TYSHtqJWF9sbn9gXWqKMI/c3OwjUPQcHn64hwD0WXqNIkcA3vUyzk5bR4UwNuQTdMR6I6k
GD6abwRLJ/qrLemzUmMayYp7As3Y9A22aCLp0DN5lPBGihN4f621r6c0PMKTnqQ9NNtw4m6k2OSb
xemm9qnVjmahntKjYurwVzibpIdyY/rLfd9slFkXjRsEnpfpH9HHOj5M2vn8zzk6RQnHVAXfgRZ8
aF9IsdDP0N/IkPD6PYEQltXk1Prxew7tTCUGTEkgt6HAzpLWmqqqE2Rs1Zatr9fnbED+XAZhg2jU
ZZRyEeJYg8Hog7DnY1OYl26MOjFno63xTLBaMHH0L3FP6HhvAE2HPXi6qAlCb+2SxIpAZmI/Yd97
Dpj8qysj+sHaNOJc/eDgVl0Q0ShM5C4Gw1m5wQDqfApH0u5E+FS6g4RLT1cwWONM8wbXUZVDUedM
eCkhblWpV4iMVJiVzsaxR5aRgYV4cSo2VWO++AYa30TUwC2Balzjg2OS9N0r322dbxWMysFOZPLG
40KlZU5qOaa8S61jqH6u+hLeV4XchGDr/kQVmioh+6jGGDkArFDz9cgx5f1ivnhrP2Jg35otX4Kl
6l8KUGbFefbSFttVvrvnYNRdkQ04p+Ui/sQ0d5q6/gxR+BlFZeAILcq1SyFQB9C/CWAM7phCtvll
IFDuVSubX/BdHHSUs92/zrkeg3NpyEfP7vk0xT+1L86L6oREpQxThHwf7OE7YZWL4yIFNXjB7w5N
elLWjR7FMoBfBDi39M+lG7Bycmp8vjUJxYQaBz6MqxJ5JCRBpSbgA4z7KXxAHjSS+Ju47+9IdYv4
aeRokHAnJ0zlGG0uCjE3NJthW19A9YVyDOiNFCoP6m3siqAhHZ7l2QbuVyY9lC6YqJn7DAjEaj3a
2/xJcMjf0rcoUcTSyCeMb+svXbOhgIXPgFtuxcS2Fz+6BzSgpA9G/zI34gZxCRgHxuaeAoW4jKMQ
CsAFs/JQJESzkVkQru9UtXgthf1wY8SEEhUOAtHD6/FmsiXUjUQ+wAXqQB6KUWsraR7LdmlrPal8
S0O7x9/2bhWWTjernyle3xMvBq46gP4FRLhNJwCwwTfAt8YoqdRfRMmgMt0g/JFh2ShW9yYfSUM/
pL4tTPStiN6qLhPKsQTUPzOv71hfAINPl0E0gHOMmbHAlnjQHyAOeUpAnrQ6pF2ZX9BijlULzSal
Qt4UkxKctUzOosiWt73xF8LSHVXy8TmzYNsMobcM9lmYYDhFL3rfSYNd0NZajqgiCdkJ04TPUXrw
qFD33q8SQuCE3o6Nd2es4SY/U4QKG/sJmQSkvfx1s/pR4xn06g8Dhpk2inI79D1E5a0GvFwfoQgF
Lk3buR4pEGD+QuJhDonVuLG5lC5YmWRKPaTcoEol+GAHRWx/BdtEK01vbT84RroUWrwCPbKQhTa4
5nayWgPPtjCRRKq0SkQmsOvrqpW2kzqIwuAKGNhESAuoEVJkJb70SddqCYeNrI7d6k0LkLL1QNE4
En4X7z6queimrnU7Jq9pjtManyo6iAxUwer1lCZbV1WA7kzXLv8k065ur8yw2EjHftM2YxawkA6t
1rOOdg0yFsthllkxoS/U9ODFAfMNmEUvmdDOarOOwiJZ3CEohDFuBfWnTZQJZsa8i0mwdYG44par
Ape0Exu7t+BO+elcpS3pEvut6br1htTZziwJa1oFBQNHbvh0yKh726R+90IXViJpDUwEAePHT/0e
+l4DFiEQkrR9a2Rc5l2ZaqKiWh4rzCUJ73tKuU7qPuEWjzB/9jm0klkx4DoL1EkzLq/Lg3WpYa+z
Mo93YRC6Vl8Jm+yUezhAYo6ftjTUHLWI37wqzD45gSVdj6QVT32xJC+9/wT1O9LqgogFj2Q0o81L
YNWaEePet+NmX6se9U8SkA3DtmALpJQWNMZjlDvLUmC5SX/16lnqfBRRkBjEB7AX7DCLfm4G60Wl
iz0sJrRx1b1Z8gqnJW1WSvQqJLXKlVJj6G9/P9PZK8LxL1L1xFj2Sqxzl7qkV/gQpB1Unngni3ao
VKzCZwhyfyNdi6FrLon6e960bGUNgNBmzNkc/yTT3DaEC90xHLjLbIv0drc5L5ceVURJDvogrFcL
ExtWgqvRTBrX7FpEXx3SptMYziP1w+L4zdUFa3PGXzwiUV4tghrFN+joEx9VP7UcmlW/b2o7pIE1
SQleRE3RgBRPQ5RjNmtiBw7eADzb6VeVu3n+f3mqW1YgP5FAkS50wrNucILXWwAE8oaXOX9pcGiw
RnOl/Hhs6fuychtPbsIRM964YWF3TCu9ftKeUxGJqXMLyyXxcZTABhNpbjc48NEUHcsglRCxd1Hw
OrFA/FUBurHKHx/+GeM6F43TzIuMa5e7PW1eA0REud2Rr15qcGF5ScrNb7S9TcXGEVsio++vwCfa
kHHrRNE6t7iHWV1ocD90H8O/Ti2Z//SSSPUXGhW8ZcdSQhQeF9ICEt2uK9YTqX8fljp0P0WrFKCo
vjaqiMjAnc8nLmowQO7LQ8Uo+HYDwQu1WzkCAgaofh3oSzWQjWBtoiRayW9zGNAHTmwxN9Kt9wro
sWq7MDT9MnhZaL5WhQWFhrLiO02boxol19DfZVJjeIydeo5rjuJg4vgErIkL1B3rKaq3m7np+suN
/v2fzSYh9Kz61zV1IhEmgX5rY277Jt5DCzwN1j4QK7tfqjCDv38I4WIV79FWI4ds195F91qP54fN
Oduryo99Y8wswaSaHUdgIo3Y6iJHtYreODZN0LBdGhQjWCM3qfz6awrIvN6x/rqIGACukiR0muGM
KXp+TdXI8O55G3Q8M8pTCPiaC09R0KNuOaGTVlLRvuec5t4mBRe4tKudljlOIGGj0aaSZJAFoqZt
dcYrBrK+u+V/gT7FjFC6eVN0Qvps+2LCbFLmYMJdI9XKjqhTqMIGHUK8T5WC1geJyIZQDgT4wC/P
swdXo+yOT5prQjig4xZlI52MWCG13n+C/Dx8PEr2xtmxC7VI6s0F0kySoEGbViWmxZxR5EbVoSfm
g9L3u+EllT23FFh3SBWJBICJl5yjAyujrxGe0E8yck/PNa14+bEVMGO73CoFwqrt3TBYIv8fdfar
1HRDw2UBedvzXXmgFmDx0xil81Ab8AUv0ELG36BRDLDB9VHEmyL7txWLuGxuTP49aG240zOjVHX9
Hv6pzZ2SzrkLm9x1Ky7BimDyj6TRLEf7u1Z4Yis+6QT7gTEJ4YpIlyvfyFalq9vKrjyHjnHPatgt
GMeNRDQhgtAfnXpgpzOLXD9Uwyzxzte0ME8c6fLcGcnL9Ec9oXXaBbSHUgrP6sn7v0fu9HDZvrWl
g9+ToThbwxNoghqL8b6YUK1oVh3SOlUfyolPo2k586tOYxQRSrohmUT45YXRFD63UDkNorDTHYVI
U4QR8WgaLsZh30Owho4eJf5njRr+4o7q03n6hwXBb9zI9ykcZZFwLABMddeZ4PKsVh43e3rd/GrW
mIh2ofsEzzdDTKNBqqwmOvpQMbQejOleKZJCPLEN4i+hLAqUdicaZk6wtO0HxZsFO/hwbHYMKewt
1IhcVFNMe+ny0hCZxzfwVg3BIVkBKuxJwgrI70w4O59UHon+Hqwu3yjX1V4ykWG7s2VsMiV0XYUQ
B51IncHIGazz4kvLTvmv9rkakGGTtO77gEklnm78vmQ/oc5v3XXQ5HjcNB1ASX8vLuSOqGH3ZCiJ
uqeNNHIber6d+V6Nq9/aIoKRSOXeIjDiNWjjfrTORyP4Si14tnCS+EOan/wlFVYpqat+nUJ2vOnh
2OOdVZoNf97WcpLMvOIqEXEdiCWGQCSicNAobWqzLVrLoE+7+efVc1l859SpwsXac3sVtiRCFLzK
7ATSe3zALxwg91LHmeOQNEzb1Tvak5ZKg0c56NvHWKGFec6ot3L4ShX2I5Lx9tyE1t5X1Nzj1GqP
sIhV3jwS7tymlTn6MNJGxoLt0+jHcbgM5+3D8AGDURmhLdmOqHicCDDkTNzWG+77KBY3wz4ns3rc
OG9miaAssuwqwikJ946AATBPUA1uMARAHsblCvfM6MvCYrrtzxw+TOU1rQ4bakxW4pDO8HjzdNws
v7kBDq5BVQ9JAqh7I6ucIqWWzyWzWjiLl9vwA4mog31Y1iLl6yun2QN8yuGfB1KC9dgTvHIEJIBH
EMQvQwUEVjInR6b/dgLCYm52+LmKu7NDugcTwB62+1PV/UYPnSNHi1M9AirQSkyTBgaUxsuv3vQ9
WjJt35/xSwjBsxChMQvXPZ3Qy5fM8elQWU6HVDEZKx2y/ePSwbJJLoCBMYctU4T+wsLmBYUJbhFz
146vtpHhSnGXp6ok5h99JfDfmgUm2uqPXV6dsyReDW9BYF+VKjQpqoSqu4KFHIdslQHv5cghIMbE
qsbjOXke7UtF7LeQDi9x0BZSvnCeJ6/ciiGliwn65qv1r1SZ0pso3ypxE2fIHgrFTvKDvK6W/m7d
M0Apt4b+rbIrG4irN4hPNDyxbGYLJUV7F5YVT8iDrr4EfATOaJ7SnzvGvV/pVgedNLON9ctl+X0z
5zgl90B6mmn+FrAEDWw63fHGE8yRr+t0eulOlMg1r6brQ/LKzD+1DIn/YfYAfHzVIp9CDdvi8evh
SMUGals1TL99cpJPURPlqpZvBOMl8C1nfquS7DpeNyVXKxORol3DPaelAdaKvt49/lAaWYpsIyLV
kzdjhTot8ZY9uTGvZMAK7hQYIzh31RKsRcyKcu2fA18/rMople7NEEFFAzRSnBN4vGWLQI9JoSm9
5alJzMm9EFK0LBEZm4EhYfcEnTa4NyqWg3+FtNYDodeQUoxqs6EUNJba/If0vFCJbVpUGzzqE254
nMtniiEyUnIcq69SHI6IYD1wz8POe+mQBqa9bvoJJyruxyEmZyO89tMz/A3AdeQe/s6ejTHoGSxn
4xUS+u7YFVLjlZqZ/KItamV49KTVQFrdcp4zDFsvABLwCyaAN1lhTchEicpbDTSPdUxX0fcnopy8
f1BWUs3v+ftbuifERK+aLMrWydwKdKKH9JGphRRNVy8ZXTcLx7FqBkvvN04qJIvyqVKfXrDjkB6d
ym4sFqDLrwZKITNrIi1Ai3gVEBDnpvjxYNLpXnBr8oB1rqlhME73qaDKZESnV1oYQl0eL9hNkagy
elZ4vCfqIqJ841vhcwHBWJ0g8KR3XZmS997/CY2BAhtEyhDgN+SY4xanQYWLpv5Cz4OIuM8u+TQD
pybvVaoeMXTC0LeCPH/tnRkgiSdHl4OfZAA1yLd3LclLS+QtDRNp/uNjQrYewcoZraf0d2OXqWsn
2iQKFHEALIY3pXPVlYwHZLkTgSHFvv/qMOpZ3jE4JKLJhUJ5REAvEEiVSNHlKyKaFx8SUaLged/l
2T4r1fz+AxAK+48EYbdlxTeEMjwHTP7J8W8evjWFSmVryqW0KhOugVmWxsHz9fzei6sknmWyXlla
HeesreUQR5x87a2Yqh13yNeStyA+BifrvOeDMTMXqen25h6FdjoJ0F85hCrK0jVrsrOjjZtIs+gp
dxdUcv6JI/dJI+y9UxRjR3EMWRPlch45jAXDdQfNaDRn8IVvR0Wfl80Reiv/XbvAE4p7nhjU0lcw
3e6Hzgxq0Jh7in68Fyzi+Mf0KezkK/O6I2X/krL8YLQBrTkTY1uSddwxd5LxfEiZjq5SYlDQg28H
sviHkEi73/d66FtZbq1Vj2AJYcPnjatp5bvmVb9L++jtjPvDqjMgNapjt1sA4HBgSMXShIslzHWO
Zu5cOMrq5IWrF52AYepIUqX3nNxgza53n9ANnc1iX5axU3HsqydBNinGUWMMkDkYl8Y3tu9FDfAt
7Fm1R0zMduqipzvOxpcDJDTcyHEqrUg4IBUjRT/s6VsBfM1IPO/EJ18eH2CF945/7pZxu94ZOQU2
RO3ICMjPBKoTOinRKafFUt6bpZJ0umT+73v7Nfp1JoSLvXPjXyOo9dLILKKLF7rmOf6Z4XK+1sws
ORrOOXYFoDrOCONOhJQLosBi8LMtAHkXXWetMLMiFy1Hp2JsRhUO/Y9pJwIfniTrMtk93AQDuknO
rYOSmrbZzmIMp5y2CqiIjgJ04nJqOCDfEAHaVIAS6B0c3dktS7IV58jP4Ev439nl7uuqIq5Tyjqs
iDcSwUoKEMEIBVLpUshQ7F+oLqHVNdpBDkFt879+GUxVnZfKRV6eAxawBEjxRjR5eCyuK9hs7xt3
zJsJL3aKBN9VFGO7bARAvt8tosxEp8nLCV1emNtMnIxLP7Pq2SADbcFj715jl21oxXpqE4ceyZcP
gHbF48Eg4Uo4dhkfL9waQf9NnyHjdVaaTZuUABXxPmm0yfhmHwTb7k/Gf8JSTxpezUIIpGmTzmxg
aXER9YCqNW9PhGfHO0UjI9guG24ZKWNcwTiRKDq/7ABF413nnEV1GzOlNHTmc2DvoT1ak1hSr1Vg
J5AMLxmBaWzFyNHTuT8QkIQ/sY1qEpRzgKruaDguvFILM16Tv6lTFvBjugNtbSv6gWULx8CNaO5C
TRL/T4taRYUPgxu/xLfRmab/lX7Zg4XLBjQ1XKYvyEK0wr4rlbhWLMT2we6GKboIi6QQBhvto4XK
qSUxeqFslM+r2RTr3UdBUjPvtdoUVd9T9vEnbwqpk8yo30X4isnCecydHTvLavHQzrraBtq3u6NF
HF+hwFTZ1p91/jUdCr4jz28onPxUUxMTnld3h7oK7AuyBxMI9Pqrj9YQ2/x/LJMBHsxwgcNss4/v
lImh79cXpIvWtkfaFqrpaYB0dk6TqbZqc4OsA3fTtPfv+kPTMe5eYgstq61RB9b1V9s4w+CeWF/O
Xtgmi/nLdoDTgDOCDAUFdvhNRLAZgaBWe/O3w7w28jAoFsy6jdR0Sdi4vzGYwrTfg1r0IVfXVW8P
aQRNjf8GhdTHj1iQCoM3zvTR65gkQ8YA0md4C6gE7v++PiAw2fEukkM1ysyfZLyi+r/fuVZGohJc
NMKgMj5I/NsIttVQXzb/NQseHH/noLq6pQpRh1XX7iehCzO7zesdOVPFL+qwSkopOFGHV1EspauR
B9P8Iv8ZPuDp7JlvkmzqKE32D/QZ2fGSocUVU+dp2e/B5M3ySBwLVnB7ExBaoXB0k9dCR2aKFFfl
8KPkUReWBLEVVtfxT89YmGANYmDPpcjqZCCILGS5TWNxEa0qz0hXh3BUbzzin10k8LzL7aGXxBS/
adzqctXzpw5h9Iy5TedNz/5MgUtLf/uzmpQjmfdt2A+iDrZs25n9/GUibOik0LJb/EqL6qtb5orR
OoVeesRqdyqGnEGsPX5/Xr5kwP7geJZrRMpGBPwl0NlS+CZCRp8FlUIKEIAlzTmP0dkbexVyFnaU
Z1uIMd7gx0UpoDEQzJYdcXEsQMp69TRhfrj88lMt+6E975NcKm9JYZ0lV0c6cVRsarSUTEakBzFH
IZlLPyxiFZYYUzSnGMm5xyCSxzZUewiL9JI9IXX8TVRCh7QJ+9qGaahV8gOA417Bej+3nzSsvEkO
QRwDsC8uJnY0fg+hghrlWcQ1eyShw+mdzjwboD5jjAnZN3+WoH58137lPRA5KiOFaanGTLN5kSRj
QMykh/nQs3xLaHQHmwIzPi0FfxAqrff2ObBkSO+x7ByTeBYE31yVuKIho7NUT7ZocmmORHWnQycr
EVJzBQRTxyfgRoaYbIHHOM/X6EjywqdHEPT8srNTW/IKu/wgzmnhECzFau0N0T4laoBpnxnK9RE/
DRzulqyEDt/phw3opJEc6y1d2yoYHJlW99zIO45BUKJcsf+cqzvTBCzHPrN1mA7897B5qFkd6Fcg
nL9h/xQqoj9YkSsgr9pXLHISUUQkm3iu+naNwIbc8slbczmxs4rtQfN3daPdgnoC3DVG6gHSsoT1
X5E/8ETuisMQIhfA7HMcFQJZs2wBFFT94C9dEC5IrhvjLuX4qfa+OlhRFXnMMG7fpnWbL4sycRZJ
a3dPyBpWr6BJlU9AuqCa3o+36xcf9vNykxG82M4veXyEkQwreMggpKBuasdRZIc+rmZVJuqs4lLN
LeUvcGLLdIgxkyo3Jt80ddHzSjC0x7MR06YjUeOKXoBTY6vhgCIZQH9YGqhGhaprIwvex6B4tLqc
CIQLedHkY6ZnaVbjxmO0jn76BVBps6T5ceAj5vq2HYdmnujdfIFKczdeMPMVf9eMVaLurf4hU+f7
7oU84fkJS8MdTEIVjoMrCWKMyRzWyK8rp+vjS99UNFIMa7RqF86Nf/F7lNHq4BKB1sxTOrvxhLqm
Z2iBoJMOkcWFnA/QtgczDkePrjezNJdZMwwbNZWttko7eQOahQDKN1NqPQ9euTeIxvHTmpoW+a1D
xsh4y7ggT5/ciqVcHoW68yLs0UlssDNgs360tvRGtU+FgKTE1sKIKjpbwr/Z+aSydGYVJ0Ji8lQU
6Hf6wJr3JzJg6L4FwWqOofXF4Qk3U3ry8FdM5p4b45dMf79cAYi2vTstE1bh4/b7zrqiCnn8Lwub
j14+A4GlrQe7jgtz7fGWHJTm3dgXuoRU12yTUouvZuQUjls6iznWjuQTOmK61bKorYkjsqD7EGGJ
BaNQvkWO71Bh4BPgs56uXwAZfrlk+IaK4L5Od8idUgxnmqRy/2RQgBeLJhnEbeMjGx18Yx91/Xsl
lVG1Hu9xQKdfTyPl36bWlZtLGB+h4InLuMNKnYgsHOF4hPf6lTjLNnLsvh6ET51Lgix12xHsFGrp
FO5ouEd0KJZ4x2g74MxHNEQcBbLkqsfQikp11aIH93d3jWsnCUwFrgIFfBIjq0X5LhtA0MdltQ/7
ld60F7SVZnCl1plTMX2amxiBW7snuLzz0cvJo+GlRHUvKrHGK0TQhUY7noW18wjo4Yu0Zim1wShi
G13DsSA9JEuFss6pJfJ7M6+fXI+pa67sGUD1FjX4fU/yVSDH2fY/8skm//7dcCJpRe/kW/0UJfC1
igVoicFvFRWoWXfpWHWFzNtdzMg0AI3324HWN/fH4DIOCwdbkZ36Fy5+ioopHNTJTfmzHNxLBx6y
FmscKknAe48CSiGP77yMWnQqT+CjbZ+r3/IAmV3oN2boK78mz9RMuHVgUrWHlSYeGov8BmN+33Cb
v4Ut34KLF1FsX27q/cBwoFtzsxBeCAciFN8WxjLOQJ8uqFBNrqcA9yaFhGi/hJA75vNaaUIuA+kp
kKALUb6JkLmZziaziMuyxboLH6eMdM7cu2iGzU1ZYx2GOo+F6+eHz4uCyzi8g711GCSGB2SYoOoT
boyu8fRiYt03XBBNlCKfVivQ+bh1DDts4dNKrwZOzLLptmGfN6A4rHmKOqpkjqUDYMP1EUlpTaWA
NNF80ez2sBVrVV5w66pzrWIe1lab8StvElzbLWKdxQcTnw3zsjNpEIOUN3sIHDb14gmftllCs35I
2rNESy/0jUJuW9phy+Kus5map2X8NkJL0hfeAmwG7VdVOJnxWUeFFwxGkhLu5Ug4eJkWwk8xyrBy
6dbebA4wA8/mkdqayHTUZoVERBpmbPhkPtVYWD/HR8+L+PxjrCDkK/gI5QVmdejhQi/mCwk2ojUz
NGV/fiON7phAPew5nJuIOaIhHiDaTc+CeUEm7nZZJUtKXNAimRTCnCUAG8k1dIglLMILE5E3LOQM
aHvOPEbSkFBvNxo8Ch2M9vbOhZa1sQS+KWLeZEDVD2L+Pgn3+HdLY+vBXuOFxfC0XSLT9HBwCoOW
I80+Hqgp1lukVEkyVVBK1lfx+Le9Tko5V5R50VMAbSFslNPjybd/ap2Vn43Q8PFu/SgwE9voxKk5
/Y/UzHRVYmRva+YNGUBMsyWU0Kyoh38b9m3948j3q908QiybQg8V2Xus3DAdPUhUlI9/n11YqxBP
6KdCV/bdtw1wX+cQhikM8wR9/35QjmvolS4oiHp/CfThlranJmArqkss25f2y9lgPJfNRmHbdNn9
DTbbQU/fMCKpTU3n4ZXub7QQFSMBGIH2CHHVcny0e40h6puMC4hKaFwHv9iHM8LaHnVRqirYQwIp
LBgB8wc+xjj90zW+/c3vxKNm+rbFsjQQlX6RR66VfQ/ZjGNBcgcmb4z94ShsQVWYLoN5OI7QDNk3
iKLp/48/Ov1TpRu0ZWCRQRv03Y3i85PKVoIserUU2zL1qmjazq2mAIoWf4CPWtJrz1NGod2SVOcO
0t5Q4ZA2787SfUmZMPtO3EI7iCVjS6Ezg2zdzZsCxdddmJwQf0OozciBQhW9QF8/BmWZVJAQi8w4
ZiCZm/qj0MO9jDtJMpLHTMee7a9Pb7RUWOh0FResDT8hD9y+Rw1efFA7tQwRtk3GdzsqTtNxRBxU
JOlgRw4WDm/UYXtKOdc75hLu1tA9wMB5589FiE/E8QIX1a1jT6R9UFAVp8iXTL5bBKoERC1Aneot
+1PTangCdmWdtS4sZ3yw2OrCOJsReRoBBO271cyowyEUGRtv78WqmA9XRqZQeUwy6g2BDdsULOVD
vuOGCDxYEkrvgEGigmZX9aZ5s8XBZanCALMiN+CswkR/499jpROIHCox1TNhIUKxoHX1Ws2VdOej
Y9OVq+JgpfSjDdFu+J422KwjCALSuKgYKA1paoWddsqITFQHOlV7dxYZNwcp54dCDE7az7P+ZsMo
aUnpCxZ/A75o5roDdsD+9y9oP4SawRxg2J9krz0EpsjHS0MTC1nAIgMH39elv1plSWSWay3DFE68
8UD/0Z8qn229RrPYQHPHz8jJy38ThFDhUA83CLdWrohzLN53s0FyNDNTDQ+0l16T/gOfkUSeza1k
PxMntmA+ySdwKC8288Sq3SDr3aYINZ06tmwxRD9c6pABd2bzxyUxMm4Jf2Ucj1i3f59rqMVMFAuL
S0D1NfITn3Zq2Yp4jKNRdFq7b8mTZDnqhXj54U2KuQDgqPQn8pMcF4XHM5zVhwdjdUXXpLXJGv88
IGWs80gamAE2eb7Zcu+20hzyvN2yBRSeelJaqMsWU9UK8Gj/AmpA/Ack67sudlmNLXOKHyOu/8eB
IrNp+Qg7NpLT0FPZUbnppRB49XC45AOAN4o2wDlFSayHb06GP6a0Dj4QpoxvHuZssGIm45jUH+ie
UWk/tMdwPvfW2VawbkHEN09oeZUSEQ6MhFv3chcPJFnqDdl/w1yKS+uzoSDDgy93FfMe/ffRWglm
0hDJGGR3cb/iCg8x91R4nq+lVCLvxreryhUuWH+hk4cREXtkE1OmAKcs9ZTUFrU/SSwqYdqFGSjj
W6E1y1SZWxfM298dGdg66owzwFldT4c0viLdQYoJMvqZcmS7tSLs3kaWYA9xdCvtuLLPSqMaly70
2+DHetszLuRN4GjjuOp+PDBdc5u3+jvtjtcSWINKq/i3wed6sg8gotT12Fn1XJ1FO+rf4oajIcLA
3OM9THv62b8/Ty906/NU/5p0TrgDN5HWmOR1EIWR5uvwQQgxKkXMZRcnxIcFqL/blB+ej0aiTRVF
1oOsRICqX4E/gZJ2ir0Zvb7UQtAFydC0im9zMBjIY4B+h8StR9ZqIbylH5kreDRKk6ohhkcMa073
N3GjRBPIZZQdvk01nlb94+RE13lRaubeAP7Ah+NZ1uW+06quVBar+hfO7hR4oHqw0cCW/oQ0EaHs
3LEqvf+REUsoaUg9GTsFZC5ylTNDUWP5SAb7d6vScuunbnqX7ZnexmSQfOW3F7J02GO9KaoX9upp
2zTTo+rjKkY8ZOCq2wKYn3qgb56iGx/sBNkQg8Q3rbOpvqg9sciK/OIgzhsvJHFqX+vQxnEKQ+jv
56LeiLURCVkL3VhUeWxE1TFUYeny/je2PCJhWD7TBsMd9vslhap+jjXF00dPB3ACsF4oLNiTG4vZ
REB9ZyP0JESc9xEO2JxO2YZnYUoHgjG9BRQpiao6pBnMhMcirDSzlVhPF4aQFffzQlWfcBdKH3wv
/IwZgEWT3yPn5jb/BKbKMlnLWcuAMlGMn5n3YPFCYoiGIfwBpocjvc+bLHALlbunS98eLPIakFsT
ULZs16MNPeS2UfW2F2OrECyxCV4raA5JmgSGPDiQ9vdIM/3ww7zeZfTaD8zTbft0U+cAbf24jTV1
9ZsJUJNuWcarlbQ1bjh+2fmBLgNjV9dfaK1WYUCkYVHz60EmxZVVoNTvdkg3BdeKNezm/xOVm69G
g0+TbemY1CFlulvM7Q9Lu5kpYo12zmG/H7RR+cxjFCd+R7Rj27SRBZ//Cet532oUF0zZeO0TdoP/
aSfXhsRRIrWIZjTcqBA0zy0jA93GHXSEAUyNsvfOGASrYq30TuDQwenEqKPyOiDoZDu95h37zen7
ZX7BTaIWGzb06yS8rT9KUnMEcax6VfVmNX7S71caSY0+n3pft+yZ2PhLdT2gJfoJdSkVz2ikWzcm
s2chBAPNJ5mp+ZkYWn6l6AAd0Ps2UYYhPTjqK79CbT7X+mdMxVoWnVB3zyLrXixBm1147fI4O0Js
pOf+nCOiEwCh5I3xtClRKuv7g2Fpy1t+3caV/P9FquOgE3tFI+RMETmn2MbE2gbyKkM8H+iJop1N
RodlaCcH9vibpYC6TaFrndD4sYpLyRgMJ1HVGT6vpv97Kitpxc6lRqH47KI+lOyz4Y2Js/8ggfz8
Ozz8EE667dqhUuiPm8wgnCYMd0t7SlnlP1kUex85/ak1BFV7hhtPcavtAXmJbTYf9/Xd6ZJ7DZP9
c7A8m/N0ZI7HpPfhuc2AFaO7xxYqUSrn49i4M0J9OjlElMUzbA9WL9JZeYUYYXRdbcSQsiR8lJrC
iQNoTGLDNOVaE+TSjAPa3ayir0y7SNEVfakA3nmjqXuG+P5a3mFplOq2EsxWBfBebKMl2N9CF2SR
doeF1K2oz7OBXl8IyF+ikzw9pq2nb96ffTxgCatI0ht5FtEYIe0res8NfLKqWUAZ+7Tq0fOsAOwY
jTWg1lAePHbHZ+TWsOy0wQu96Nuny2pu0gBOsi/osGlDoerb+TqmDxwqD/kwIeXMDVoEW45D7onk
8qqIuhjWpDPs8CZzpgAI0uVuJhLL6olbxLTMY5ACnn/RukRgeNR2vxGwCip8VA7/kL5QzJCz8sie
nGG3/B74A+hOQq/QXIu9yUM0OjGkhJ+AoSqKgc+D9rrph1yFcgjscnq9QRDM0LAdIfuEfogpv8UR
u/AL0mbpnRX9NzUmGcW5ENejwUchZK3ykTOHfdtfd//yzsPaImNzgNi6KCS6uA+Z0xlDcsy1nGCU
uALrj3CZ88F5EfXTLjGYDyaeDkeZrNarID1hLwuQbmsx78PeIhY85688O93pScMyLnPnBz1y4KaA
pN/Qx4XyADmghl1xz6KGfLA5mxGKvJcIhSov95vpn5tVHtvLRrEVlmzNssrPcX6bE4yOhXFUY0CC
JD6KpWBM8jSJ24lKkrZtJqY3T0ytz89cLwhNuNr35tNP9ewSNoDwPLWfmCII9qfVRE/Qgv0Ht6eA
5Lmq+uG/hei9fcRd5mE6buh/24K+FCvZHv4SpxNxx5Mly090MCxT4vQqRt7x1o2cRGf2FKsbMquf
/358xGc+0UvdPjmWOD5RlZtG7eEzwp7OmLa7XI3Xd2RWA2zAZ0pHWZhwZjow9TTDPscxdpllLZWH
g1kctjBP+4wwv4580tGxkj3pCGV3GD5L06p3hQtk5WMFis3I/qYAlQWoQBi8gEzaxWdmAUf/5rKl
RREnOFgdvXBU7hlf8gjhWXdfznmpli5SeChBuTRW858ghhCh/GIRFP5sWaeLIhnHwknGBB9cFuzd
iyhvWJZYqXZZk5WiShCjhJTawnG1s5RzANsdIe8edbOhh28cRFbnF6ffdLPxl02yj+/tFFmPCNSI
KjY5JdK0pq/waocN89UVn40zaK85/fS1Q1QI8ztQDsndTx2U8XnsN+aOzODZO8bbKkU5zof9cuZ/
ayWwa/i0d2wnXvRr/RjwvcA120xwp2pMdkUkx7B76fAh++dIQweIqd29RUpvseRb5apQI0ZSfIke
S7BBunfAcyjdoqZQFLsQZlnR9yLc1lfGjHO9wz9xfm0kL9jrG4Q7zzIir8+MWbHfJzrC1e9jE5JB
uwMQ4QYqsVL0O595aKJvLCzitueIBn7ZoGfsdxWWC7sXhSFSz8brXQBh6RCPXgURuXWdDaBV5cUb
Q2OE0ldV6bKuW+H47ulIDPNBK0x4ZJ1SqRmxxJun8I0+MjfyX5Bh4LG52mXvdiAYAFSNRDu02itz
9O6Q/17B+taiSRYZoSp9AZQT9cCSeEzgaFHJT9yR3WI0Vj4Jja0BWByx51noUqyS1GkMAkFf1QXe
Ne2yJlYbxU9PKwXrVfDs9eXke3L7+8q/CVYa0qLX+f4pjkWhZM7czRkkQ9SlCd+aKf7y6cZhFPoI
a8Bpk9rtCLYd7Wh0mZB5h+AqJMaJlGJeImiNIYUwT/FtL3YYRWygCF/CBDewPl7mYkTMxE7JGRXP
68czaUExc5EDvb9qLzPoQFl0KqqO9qf1lMKWuuK9/SrwfufeevDYxwV3tgbNiqKrmTy4xHlJIIt4
hbEhAus0g+8sjGcXbRrX0Fav8EFEeRK67PlAFgjqYCcPyin/SeMRr+Vgdn9zalzGZptYH2fLhDeD
n4/jTtFO/yeg6w3oR8AOg2yl5gwdEVh8HfhPXQRTtxt6/zsX5e9tqMOak4vKTG33ZoDFqmohPvdH
QGxWuy67Km34YdPTUZqYP0p1TLxnbtVlGM23Y564sAh72N1WNreEU+8todwT8PrULFVjgviwYI1P
yD/DOQ16E7dIE+wYXlr1ZBrmB2qohj7RKlsSmmOy5PuPVFnlo5E6Z3DemiR+EFohFJ92oxQvntCy
oNrZzhTtGpcRb8bMVEpmpiEbwyF54YcX7TrLgzrtCemd6SbeEdcw/8q1TWkWTZOOVLCq+3ExZLnT
fdFEWPLdtOjguFnQJHED3sEJNb64g5tBEW/jowcvz2yMTQqZhIyDhInXz6FGZrDUPTna8j6wpOY3
vAmbzjbZubBDPd35CNx0+SiNWScb/xGRkou9gcGmSS0H/ZkWrVYGmetZGpVEz65zZVKI7IsVkPAc
qVCuaXUx/71F11zjRR0Q8qOSRGv4EDKLdXzwx3CjmdFrglBqk35Bi3wQmfZ3zRMEApY26sAMmZrY
K8PbLwdN9xirOKY67erCN+fz/UQgZg43WqYTZaqsY8orCl2c2aRD2melKYYVpXF1rGvzOAThPkud
ucojWqxc59NKFdVeUjGBG9p95hCyyyRzYxZvbJylVcKjvCQaa211wgHQ75gh/O1tH8O6a2hd62tf
NjSze/FDL6athCP9/yeIYQeYIdIT7Zr+TENCn15eC/U4s71f5sCx0+wLXZidzPgzN//KAfqKu+5l
9dW50cba7045cghzJpW1VtQApxlMwxDTzBV/pITC6Jme3lf5QGrvYycsBUA6LfxiO/Ov4PaWXrFz
af2AsGsnmpuWQSkpC6P+/8PRSWGVBVL6Oi4MO+uJY7qcg7JLetDPHiUg6ErXp0oCui9Trz2c45QZ
lGJRZVJ+5sOSUkp/qeoLpjeJo3/bCptO1ibG+ARxbRb8ym3/0wyw3nt3/yVsjBc6aP9leYyttxs0
bKOqtij8coa8DumTrBfKQespqEReZq+Ikp9pfdl/qpIGNqLxsRlsMCI8KYPxcqx5wNSayJf+JA2L
6MA7ChGhIqyeOkD3bByjzLcvGicSam3RkbkWWeT02bU+t/5PwAKMRFyqZ6SSI0u8rMI0sTIgWoRi
bZdcpOxBlqEeVQoHHWxxE6hUBdrE+lUFJ1jFnvhrN9nN2bMW0389ydi6MDLs7ZmBEddQUsctU7Ri
ytXyfiDZ+HUMAAduvaQpr3y/0AFw4PrriGorMrisyElPoMjRb5dZ+bl6WVBJqRKlb+v16Ya4l9zr
I0Ni64tGte/zspavfxwpq+Z+dNSwvVKkHoOLZqO2wM8vQQPyy2GgwMC6fJM0uib4aGrNDT5ABezC
0v36qKNz46O4JUn17B6wQ7Gf9Xvf5pN/sVAknQ/IebGI4lG4LLA/1C9asUSKMf7mZuFz8UbNSdcV
/vn6tkwPEIUnAMQUKrom9rt7ujo1ekGSiqqASqAPJ+VgoYRLsBNIBLyTj3srSYCh+diCrfVC1eUX
7Zl+huUbMVI9MPBX1AeA0fiKEx6Fy68WOJkA5KDDbWAYDnrnYAcFUEDRdR0S45Niojmv5xllxw6C
9J8WWHCtbrgb7VLMqQUS2lzzBU6uC+b56ZWM2PuWicPYzg4xd3pvc+1dRWgK4CXeoXMbjrl2idti
Bkl9+bBko6Pgi4u/aq3AL181AyXxhkigCmAq+PgEHQY/vkz0aCkYK5zu5sPZmVNPpdaCfQmaLnCA
j5kxrVNM63hEnj5m3PpbJUOO5gRb0h6znivkG7MvCvl+fYeCcBjlFowlkfAPJbNFiQBqvsZBhG/K
d3thcYaWzj3a8yhLdluOuGqwNgSKCmc3Trb0nOW3isDKmQp4epuz+rAJk6v/a07e3ypCDXKKGb4k
tt7IjJZOP++6ZuHDYLXzx1RzpvrZY+r+0WdMqX5jTUY1CZ8JmS1PI8KHBU0WTIZzDLTTvYg4kul9
tAjn64ZxfcDQrO55ZL4aJQfd1Ui44eUtyzv0JfynAisKsVL9q7JCyd8M3sTGx/EEedQAhvE8JAFi
XiGbipuCWYO2vcfqSm3NZPXUGVbXIKpIK9LjFh6zwJT7THL5UUYQdFaURyqSdw9OGSuEaq2giNh5
65Egkrnmz9KUwVHzvEJTFitb2YDiItFq/FQuqyoH5MvdjowYp1UONyuq4tVT4rBErzLHQwiKwH2Z
+sxiq3u+5NbuNxSZ3BWsQp681crxjDtOxmcqut6+EIwInu3P6b/+EVlytQg0fvXSScGC0i7aTtHm
IiyGgC7MnXVsfJ935+NeUTBjIuRWRqRqRImi5ERoZgYb2BxxdIqMnGHgcQ40Xb9HuZfyU+XFKPlz
56R8HqyFo/3xNbnKSPFGq/q3eyDXmTgG45qK4vSNKyQt/cTPwjakTX9S1tRxdEN43RbE7hRqScDS
JF5UN/HzCmkjFNQoH92Kk5Ij14i23m+SdR557N2HRvYRB/3y2b0OXph4Ynle8yHl4Ib3AO7U+Rqd
CQ416kHwXf+A2RvSoQG7AtHAu876D+UhfGD2YhCp9Zg1wAtstFpUvEVbl6wkzrLoN2LgwfHBGA05
mvsgNNAQ6+FaLyfRmODwcXuAceI3iVtpvFPr3EQ8kg2ga0RydKz7qJ2FotAkX/3SEp0DG+KMWvSt
M13aryYV6QvYyq7bFXtJzc6b58fT4ZIKrAB1BlC76cbCXOb6UwIUAxGq21CqH+bWpq1NVbM/8iZL
7vDTypkyGn/sLdASNirRbDoPqbHDqom+uiPpaM4HICsqGN7Wb0fP9RaKYINmw2h7UwPVWyssux6S
5mbOiDnrz4jiebJJ1991jt1IHTEf7Ia6nxcbOxVKBG/GYcldrZeZvUV5IVktIEIrEK5BgfYiZeZq
TrkFSV1Qhy0hspTBERUH19pYlplts5G4JADQAevjjGP0eFvkp3pWI6UhgiVDzQmzNw3DhynSRKCr
fhAj4xh6p7qk2hxwWHrF5sqT8cHUk8F43qc2hSDgEOZtD2u/gcZR5wlCAedO/ZblFePJzNUDygcn
Tz8R8i3UUgzGTW2z8Ge4OWQ0DyWTyzd3BCIQR5xRxQydAj3TOvSX12x4wLk0rriJo3YHqHZDGWZw
jIigFDfurOKtslbVrsmJDcZUceXBc00121pqTDuq1qSIA8KVTeOivPAqyRUT6Z4fOawb/hhiYRRh
bGop7/tPaDRgnHgRCvJdzxteHBvbGognsk6qJ1mCN8ax8Kbw5KpdCMkV0qyCVToC7Qq8F4Jqu9J+
Nj0b9UAV1C8e3QCFA27zxxoc8UzjzSHk8VxoYe8OsY994Zt5RlJQ5l+6FUYmD5zf2EqzPJZ1hpDh
UVlZPq7jQ6JdlkmyF+3Dk2OA7CgsbW2hTogbxvtuEWKeMz6B/XGJNr8+gILrHiXYTz+C9HZSjRWV
yIym3d1oCTRvt93tFBwOo96DPIxjhMWQLeSH8KJh1lppOZtAFagWAmu02M8HGzzui16/bFP0ryWT
8FUTdcwvnBtdjZP7wRUhw46c33QpLz5AH2NI3ZzSXXz6+B8Vov5bTbSJt8gTXqi7lTp4kuSUlEoo
JcU/UXpqdCkXZt4LdwmDitNNvDTZsiaLaLQ95tIcZ5vo2TYNAK/YvYBS+kLgpcTxHMV+srAyWSOk
KOpSdEI3SaS6O3I23BLzcu3V/4EibtkYxMvPN5Q7vgANwSNbV5xUiwqyQCkr0LFVabrrvFOAregI
PVCiWufFcFPjArmP5iU+lZskGABPXvk4EltnEnwm4DAum4ETXhAD4hdj6c7bwjq4vC8FcCUWjtkl
TRTFad2iUntVtArJQd0CEXGHXojyiRsIb4lm9r9cOI7o8sbLNgvQpY7SfnvO2BkpLfp44iBYHpB0
Dp1eXd7VpEOH6pokPVvzJ4m7/i2ABEZF9piumOO5iD9+CH2iu4MYaOph7pO96OZHmZDuP+qUmOK2
sdI8Nju209mf8GpGdZIwfrlyjnkBZePwait0PsQlk+ZBAU9jH2BVibSjWn7zuOmy3FBiA8udmP2/
wMVYz5f9mlZAdwT5FywlW5a0O4xBiY25LZWJnM6Z8sC6MmvOesqfR7Ze//VQvn3JKeF+Rfzmb+DW
j+GYJ3SDCsllXfRjieDffDzJA0g3Dk2Sxwlg19vUpcaU4NqGLNjjzVuq4wD+v22GqB32Kmuggjh9
SF3GYEaz+wkbBvzsbrARdif/5ci47T2WRfWhoUEMQH13e7ObyReedq8zAjVTULItPvBKNeZbD8+o
60FLc8U4V8w1G+9jw+0gUfkSpVkvwgRkfb0hnb3zHD1FmlEU6+UNq8d138kZcHOdpgPlfW5sscj+
+USl//Wcb2CLVXstqcU3kG/DIcBd/A6xh6hUHvMaO444UbrpIOAZcT8NHY/m8LyaxxhlAM5lSFIc
5n6wnMPc/NW51bb/dS9rgsJTSevsxPmK0f9zI14tULiA8YCbClbVtc6qUPKOkhFQ4pDhAc+IV+K/
5kNMDcz7lQ5/7JnwuGSWBBGeEwqVsMnT3uKXUdyUhEpKfg5Q31lvKmAb0n+lTD3NzMgJ8hSTiRw0
4n3YBr9ozw983awkpydgqS72tomN5xh+STno4mBQLtvnNDXQq3vWQHltnfBoqZeDQfkrL6oHvaFn
9YHRpnG7IzG7jMTBn2ADAWARRzxAdXhDtzCyP8SmsaMFxwuyMKmr3/ezwJdq8cuS6k3+H4/vn4zQ
m7ty5EoGYSBf0QI6K5CpyBwpvXUpxV2n/XSDhe38jIC+r9UR4eZreot//NCcJSlwJhNiMcrd8e6B
WCb6uBw/thDVZ1mnQ31lbkEs2IQgMVjpIM1blBU7HmaQpa8uLi1j+8kkXZU3dHRu2JfhN1jxO8TH
5p0slQ6yu4GOs7VJtEmRTQKAVzWjwL3Z+C2qFLCId1YUvrtlPfFpBZ6KMFmdyJpwCljQDiTm71uo
2kKjpjKOc9DaiATImFx0/jn874NhSu4wtSFIQsZdxZq38tLMwMXyjOPGo3vP+d6Cj6hyzTbqaKNR
OURQYLWHf2UpOoDt878yl4rH1flyLL1/w3zsjaOX7EzFL7q4A7Saf4JevCD6OOjpCRDGIgZ1S54X
v6cdK94DC2J8zXw6v9Hz0iv08Pl2+4KUsujblLqaIFJnH3YGucyZ+r8DaC2GwYKT12v/lpDlpsME
oPxy2YhugP6DYBjtUsdjOpQe3PTZ5GKNOtHSpLDeW2+H3ZujqdC3ZDnKAJxP92UcyjPXcDcBdRJM
QOZVkQokcFFiHl4R0o632NCYZSVeMwR4fh0/LPAgZPR18+xy2BSL8L8pG5SUZHhbdq+plZNB1Rxa
SDn4feAUlIGIdvpWQNiLBdsHEx+NOvNCD7OUduTe4tc6gMmLsoi+OVB6V95vOAYPbeTw42/KJfHK
KqhJFI1dBcNdDO0xxbRrpKLq6plj1cAzOGqCfLRwEy2yyoTqmWGxrKEdOTRwoFbi1FYSjokeD+Ga
aZcJAXIHpSoZdMKMK4lSvXr3micBtjMytOKDnuwqsbpdy/740LyIYqKp4tFMTbGNR2Gz9p07LxfI
vAPA9ZhNJk9XPL+X8lfKivg2TvRJJozxNfA7MTrCiJsEZMDCoRavQT5LDmUhSwEL6NL3hGIDVdr5
qanhELyeTGPxzx05prfeHHzf0ysdIP2uia1OyxtZ5hkA+FwdGf2JAj+1cacZQ6FPs7J9hEAZ5Ch2
WXuC6Rmg89JaW7YosgX156We4aFphl0MxGgww4/YunO/UdlOSb+66e0JS3ZbIRCWQwtGtnX+gd1x
P/7wCXkouenRvxj8P+DbFIvYxaQ5o8lLDA0qFaCGxFo3Zo7Kch4bASrQSFyS3ITz4ZAvhqmhzv8e
Vzf9pVcP048AN9zXkQ627XlmHEXpZNPzmxBygRd3O6371f+ue7zKB5oQABvrQOko/6WNJfYZl8+P
k+pSHhU9cGYof/GTmjKVnJDxvhtj68XnV5tNVwst9qy4FdjNfLCDjtmNkQAnO1NX4T5hQYfS/Sm1
+uTDpd7Ds2lALR4PaLXMWz6FMvFcignVoXOnmAqfGaZ8mxZiGpzPmd7fcyDlyH4UXmmhs1+1iYZ1
FRMsO4NvfKfki6tbMMV77KTcb/0i0COBzhHCPI6nQqF9J0/86Cqq9AXmqRfybu6yYRM0FT4UBaM0
ijPbEaVaxnE3+VgZgE62xNDKRokaVzDidTcLSPLP3chZDxb9wZ4APr6kTCvYdU5Ns/mKyu6OAWmI
Ul7uNV9hkcLMONgcYCb0AU7RndvXRK2ktxs/tcrEH22xVyOatND6rXm7FaBIl6sV+FdDJ0Nv9Z36
Zb1kxXKPU38LxF5CFwfgoBTduPrKhRPoN2cjDsxfBiGSuyLhkXMxNO1CGbwJ2g9xZaPtUfdAZuOS
iSipRxtcXA3bngW5EJ4qFYwLetEwXFwoOnK1Ri7hNK1VMinP8WcF8NTstNW/mMjabjJ74IOpS38I
jFIyn++kTZZNddimbRANPCTc+dHODX7css4jxtFB9YXChGoMn/MZ9Jl5SjHZmZQRfTUSRNh2T9jE
JmWZ3FHdoPdMZCJ20SvpOTq4zN5DbuodNl856qRwXA98blUj37Sd7OyMMksnGFUYxXWy4Osqy2t7
Xp7H8fUlz7F0xRkPjGW0/jGtau5PJVXOg/Lrfp0fmq7D0hVi97Ck4XazyB70VI07pXGl50CHHiZk
T+E3nv/7oX6KGi5Dr4pTcFcD07HoesoWrFiJbhHlrLqsIdCPa8YJFpsMGKuoJlu9fLQEFSWKY5Up
25pt5PydGcitx+C5POE0SSiFKgWIuxasQNwKbBBNmlZpCsihtNXi4L4pywRtObJ/todSEiIryiOM
A4gMNWiVjUn4SpNmalXwdpfQqvBHwV6c2eZVBxWjqbFmzC43HnFXuvRWP+siMsd6qViNIgRM59YH
E6BNNAkKXupLx96LtZpdEobbCNuh/0a4JDLMd2aytHpL35jZI5gFd6dSR3+reTidwDui3qKxq8+S
QxxrcQKBkscPGVOSfoDwP+Pvbl+YDEmIzZa/qVWbQ2dKNtvRVKlmAh/1TTOxDOKpu9M8JdDbn+9r
PjHS7PjfrlN9luNqCZ6vVHmO0DKwr7rSz05tCIdTHguxRIek2Ozx0sgIL0d+2V8a2vANoO+kL2OQ
8zTfAEgwV8AGJMR+xgkiRBvaZoxVQ3Byr3/NH01aQr0H2SWTGiwS+XyiZrrKwdqpsKXR06dr95hx
HkI+BmRIpOlCPwz8owDwsx3sJbpKuiu8IVYQAAOaO8IfX1THgmhGIfaAmz5c1J52r5PbY5v8OiyI
kEIc/qKJ4oyQ6PYxobMDGV9OKbq7Q5ZXqfkI/k0C7fOOsANZ4RBbTDWhr6NMB+Q1/E/tA8/RnFpt
2qkvI62zoi5aZg4V4/OGz5NdQfPiwhVcRRiHcw0/jNGge9lw+9mI2RpjNyuBoI8yvl9ecogzX5pY
BSk9JafwLWZ1tBJhjZ9k8q0hWL5uzHSNUn1LJHIcjk/LLk7QoFaY93/AE3rMbxtsWILoiV07KDwd
uSfKZX1JkJK11upMTF+KNhAGpg6vsW3NKTQn04vf1y47wC6Adz61jMGF3iJwQED8Fk/+zCnRA5Mh
BQvYtx2GTSb+cuu2fkJ7mA6G/xZbKiIdlMuV15Iop5PICaQcqq7VOllP/h8vm6dOvsngcyXmUnG1
bnnWD8kKCD3n0buT2RzzcZa9P6PTQ6K0UtYjIt0bwJou0rYfYHkio3h7D6WMC+XJQFCRhAMpnkvZ
t8XfCBdoS5eiekUHTPG3O/uM8jvaie1ge1wyYCa7jZkGy/+tZO25sixw3YfRjFOjnN2GNeAC3mtK
7FiNLmDTgQrVPogg4bt9IpxX4MLMJ9gK8xVWCiwFRRlYGOIi56hMMDkYPKXRhGRG1ExUu6BfOfy+
rXyPzYx0ZUqpzvXPgQuIk07EWH7ZI1sdA/w6nAITW+DCGHYKD3h05fXCsxBtf3xceu9N3JzsRYb4
0HQbcDmOpDopoZ9/eMoD5mvVyYlw1d6xOiBDLD/eGXABXYv5ng0kRnEFFP6grPgYwfzQ3T9pKSUh
oenRujUa4C+uO56hb4YwRkXS/HoGklwb2fg62CjVk/UrJFGEOLsv+FTSJ9p6hjpK6xCRvFhxTbFc
6F/0CtKig2vhKJwRg7jBhhhDOJyHFnmW9Qcwau41D59H2BSdK47PFnthyYbE66UnR+5Jv4deMuwl
Ze3YUbWmJmrCStqHoTN5EQ6XgKUe7NOXvqtZtBZZ+A6uijLK+okp0SwDhU7KWgDwwyH+EOo7NGsy
wCfkCpMlIaFVySTdNgEXel2Ykz0M8uA+6FyrpmUqap9AxEzXiR6R1EVFxo8V7SPqwSLe9ew0TPdB
hTc24Jy+DzHXBrz8RKOt81gYOLawyDVET9j7fEWW/gR3/lsIuRICi6irc0cVd+eXu8LAbtCVSCUT
FvAxsqWrQDkln0kxh0YhMXF3fN+28eD6M44e36VgRZrxRUIu9AWh/0VcbVYxLjtCK+HJ94lbRNIv
hRB8hUptDD+L/62ywYtLkMW04akyFaJlop1rH0LlvhlpDz2CXP09h5JKyrnUbwUVo5sJ6WsIsk7t
Bqow5GduCcPvbb/EV7F+CBwPkdX/525voQeln+KWm0j+g9/Cti7x9sjERfWKeTmEckWyQ9C0xDfN
WTiH3VCxE2v1KV13ceKyYTsEFVc1irUTZKIimlorIPye0JytKinnTHU8/3Z5lrHzmMfpiGcuwxgi
UYRwlptMpUu2t02GtKIOqzGoIo4MezoM4CounXIgIRvZrudF8zCDGQIY8Z3kPRj0H4RrQXmK9BP4
OvyihDa0rO9yOO3Plf2hThHPZ3hdO7QLHgAoLZDVu3LvQCqzCKxmM+yJ3iC+Vu1r8alluffa4YGp
e0hsMzmR5tFDXqfQ3QR1CXhn6ZIhp1+09T8FWpOom2A7VcXNfjx5dcPcpwvImop/Q17xRL6wQKFj
MsAKi5T2BhbCoRJe9+KZ84nukummyl6D7d1hNc8oHp9ZrJ8YchP4YjPi3+j5icDpkkAtVrULzd0E
KxEv2kvwid1DO+7Nd/G58DA64LM5TCHkPijd1MHgx4iUoIHqmpDVUcLHGu71VobhGVY3g/ENTgIa
oujla9BRsjmCvum9rHFB67zJSA7JSKfc7aQKeABAAxU8D9QeVZRE+/vBPao8b7mrxDxn71dgopD6
+xHRyHuJ5h9Bl2UwgvzMBrlg4gSeIbjM1zfO/ulzwjx+pmVbZk4Kaeuz3L3Frrj5RjG2eUe+jNJr
9odICxAEK5Qoe/RFXUFbvWWetJpUymaNUizdQp50LcJoa010w4Tv/lbHof5o5IIWu2ZIL/x7LV/6
FJcfNuw+BYlX36FYs0+49HwPKH/UsLQiV6ENjwjv6W2tSwR00FboyWbVBvUSqoTNA8Ikz9LN35iP
d+01Gn7pUnt/A8fJXWE47WWjCeK/r7FnXpSZynUOeUU/Rb1nc/Rzejo4gXPKbxVYDN2dJ4C/CFiL
Yc41hCxysub5tKRwfoIVlt2ZGyyAHAfwo5tIt30trlxNN9m1G6FOK8eEgkQF0z+/MLjcBd6Ggqoj
vpG1rZfuMqxIUrfzt7BDAtV6Km2qVTZ821rpRasTNG+SS/XccvXi2ReW/ytfF+aWXBw8XueOzQC4
MHIvz3DegD3WLVFvaQrCUTSET97cVUyfa7FRJmiDaKwmJbIc3R+dLrNAyHhjIOoM8UJ/RNFhlxi/
AAyBPzap+L20gLDDtpwQ2Y4iPTDStLcDyQ5S9ZV/EI+V3ehLKQiXhxUp26iXNbGBqzFFwf7ULPn4
82vBBEBPTGvTsAl0lj2RxJKc6bd6FQHgYW6woiv0QkmTiEbEFj2dBLDJYEUenBpYEcezWOF9wsup
DPOr5dtNH27XUTeSI0ZNe/gKF32VAn7pkHJ63ZeWn0YqvZe1L+7BIFLXICQXrZtx5V/tMyoE/X6W
cgZ1m1HWF64uVQiZSDoe99ROfTglvztrx1uCVQIHwXILvB+ctADBoloPqtWr9dQvqodIjfhmMXJn
OSTcpa7tLNdzgAx4bDmCYWKhlRmIzr7x6+rYpq1YgJduAJKYjD0mIlB8JEXqFP7eaj0tLSlFU6iR
fMgql0ywscA0T13eJvsw84eHbzs/Hwg9QX4o1A3D4uMK7oiB+0+e7eX9iQopy9keT5SReRnDU+dw
axD6tGO/ub66q2mHgu9JQVg7dflRlDqLfJk6opRWikruO8tRMD0QZhngY/l6ozayd2oTV+GbrwFy
slTnGBcS2IN6eeh7WQf+oKHpWclcv47q3iKWqjB3Bp4Gh/E/DHhGr7WcMe779ZCSqyobAXAQQlLV
b2Hiig8yd7OPYgt/wOr1doS+Djn9X5dND7P0oANa86+WhpvLvwJiDOPgoDyGTm5DSIvZ+Bi3Thjx
1twTdBad1SQ+UL4/WKmYRH0o466x/3n9VCwlRWkowTwpux5jAFcGeUOr2ndT0Xi+Urk9fbyQ/Phy
ev+MFeTJiydc8g+S0NmFs6C4tOTbyyodM8YGGVATTyKadFfq8EAD1pNTmkIjBI9x6Q3JpTd8N72d
gkfwdYD/3WsVGW3Q3E2WpgiKvzZ7n9EGMzzlbcvhSGYmMswHYVq8k6MrdxysbvYtMQk6CRfIZ/4B
ptC1NvOMAAIam35fEgrEA4edo2wiq9iiobaSYdQBnS89kTLLxtAhIJo450L7woUCj+tNlAlDr9PO
0oTHJQ0mEpP5EDox0S0HLVG13XpqJ3n9YeBzCRenE5+3LsVJG1BmcriFYNy3lwJCXC4kZoooHdCr
sFD10LBBiRKbf1nXxo6hoB1bZomQ09OuDbfJi0sQLzcxvx9ZUr/p6WaUdNBYzLsJhIZpUDLgVACv
t5c93ccKKcvlGBHj1kdQ+gJwOFfLFtOMadUJ/gv3l/8PQW3wn+guzgTG0OZwNerJ4NSmgq3IYk73
3h64OIAO3xhNyA3b2gHjqlJkOi0u47+mU8l8CXjm4J7ZoHcpur8/CoCnMK9ZtfXc+GL9PV6PzBJP
u6Ii9WNrh9+yGWVFxlSmlRIyylt5okyUcxJZuN69hHLv5H66u6/BLqnJmflJXmefn4+5BSrLKKl3
yPS+EX64JteEbnrvcgFWfxO/9ryN2HWty0Bi50BJEyD6lZNUWOP6j0U9UzMcq7J2mAR4hh/ojiHE
/9+wETJnR4Sai9LB3gbGGJ56vL9UfD7eAd55rdB6F9g8Unx/AK7PP+vpTJhqG5QDJUKgq/W3t1Gd
+NGMFbfkNOeh2XPilqVrN6kEIoCZ4xQDzXbZBSK4wzOjiumzC4Xdnp6imfjcmLvGxOyB76yis6PA
XfI7rdl/f7CTAENENI1DDq5dvZA6+vGHcEdHze0iXaXEMc4v8RVYVHPQI4L7Q2w+ZiWEmw2+A1wE
njlIPnmXei5a5qPZfOVxe78x7vQ76J66hdeSWI54ERMNwHcIx9LRUbuyQliPQHZygBqWua3TGh03
NIXgthR8iz29YDj4LnkIATeEYKQiD3scw7fGDstXFH+J8YChlRSmSVa/uZ6hFrCK8qgNdZtR8ENv
eWAkXKM/sTZYBYdFj09f4JKAwj+dxVM0WFq9Zkx/hUIyMk/c7BeEfcxRf/zjsnYP28Q0ZmZH+2+A
DN0klzBELna4HqFnNDMAxGrl2dYAysFeOLKpcnNLfPPU9dmjnY1n+lmNADowrA3oEPM8IhdxURdy
BTcG4Zow2Tcctju92fYKJf2u/0XknyaMgWh2fxhDlVnkocZkbWFonaBgMRVuwzKWzBcgLna813lo
R2/09epqNfSTy/jZf/N/cot2tkdRxK7v8GPDlX1FQqnrP6Bt6P2xLVf5IeRizX0xtz2jy2H/xfHe
Ii9U1qUlWLv+UL9H/JjlwqS5qqS5/NjIt41+CcheNdGUktxieftgAcDD0CMuueHaebpkxkA9Vsou
W4v60SiMXxLhQ7AT/zi1Bv1Fvd1bU5LkcSvcjt0vPZz+tDNOdXufbXco4jIkr13v5NgYjOHybr/H
iePGjI7BQiFac/BchzLVE8uVIERH41dLm8ZrwEJCEwcYmZb0ROU0ufLpjap9CXlmxmzu98D9gSJm
KpWk01asEIS2QuydbHV/Ye/lN1MIAPQp0H1ZTgX93qK+g34S1nKZ4vdFYSxnfax3fAuuReXOGcQ9
E7rOYOqSvol4FXMVzmpCOAgASrfNEV/4ilnBNMup+P/gh38aNBaS0UrS0+YiYWqEB97k/qyUemqi
Tjoch0411P+ZOkmAR9m9QECmtHcMlyoLCe5uZUIYzjq7jjGFS1IJ6d42oevfPLEmxeCTBHGUkHvs
2m9HFZfl/JHjFnlAIspCGR/rVcKjSZIqza6VDl6cVpiOP1wenaWjgPQ3D6Eghk09Xtk+3jL1p2CY
K5MDY/XLTHxTAG71RpcgIliAxK8SmubFnRV2U/U0gXitYLxqDz2oXlRBf3lYlro/VFL8kGB9H8ni
6yrE3mCmNmRJgHEAVGQV1S6YUQ6Uu0QcEgNOVDF7oklOmFp2iZtEPTNbk1Vz0zEs8gDDRbvfsdrI
FKI++MhIVXOHtkT++dbr1cA3zn799TC6rgwwat7vPnfmCrNI7Tl+MphqzrJnVfZTqTFrcNjCblb8
0GYBr0iQUyd5t0BrKRzjQ6n+EsNlBDvovcCtI0iNy/ewsQM0LXB5kM3/iSmfb5/rhENf/u0bpjBs
ccutGbU7eFtGKyiODVXoSCh9q/bUzlrwedQN4NB+iOXhmuF7XYGf4aJzZYB74PTxeAimTu+leIUb
5N2ydFPXiWScHG/UL97pj6kMJcTq5AoxSZzy4g7BSEXqVYt6G6S7HgS/Yn4Cxx/haNjAfsArDZi/
VgmUDhGzJQYL7qfOj064EqRSkir5gArwPVtStIktmOzQI99EmaGSMsAS4cWFLvtccnkeRPdy637a
+RI8ysVG0HEo8U/I0MjTqaHuOSmIS5o2kBWg0twV+JeBQMeT1Cqm/8/jd5tamBUvkninG30AgDlj
S+PfW6/e/I5Vr1eMzxrHlW2kGhHRvNycUHacT8mJCrU3Y/UDwW2DYRM4vANvUYDjKPxtSutDFBJY
dE1GsJxlRmdWIWh5zfEYdLMA6xpslV+OjEZS4DwWtoOO6VHRubAR2Ofpfo1XyUPOVrLvC7upIrdX
WFNDVree7DVr5Zebg4/hSWLKA61eRh4pH1KEY04sLTRKJIAuZkHu+YzueAmslzWQaCTRQxyzqL1H
gJbbe0z8xdbYcqruX6Qr9RZjJ2KHKQv+ugwClsXx67ClS0lTzdLNGzG/Ga7Ig7l4Vgrak6ZX4OsM
4VMxbwDjZq6a5vB834KcFviZpU16NdupCEHxE+L8IErOKWSO4MrgnFgN8IpfeSdPSy6Jyp5P7Ecd
3JrGTqw5JHGyK0qoaZS9tGcaDcnkZXzdom6Hut1lcgcSSV9IZ1boqX4mB4DkYi9TZkcIAgldqdLN
+OJljgVprms9ypPWAtrVUTMGLjSWxM+bs8kXme/h/7mBoycNqu7N3RAl4tLx4gotJZs+YGSDCone
4tzASuBvjUrVM52OCykE31ZE/Ng9F2/mVNyqo7aW9w90FSewcjhqIYS2w6fq/GNPgsV6NM4IylSl
K4nfdRFrr+Fg/B4oXFIMt6BkOwVKJsLBsR8FrluGHhqCXGdE0YRk1ua6p4d51ce/AG0n6Tg57kl2
bPmSC+e3wknBH6h00dWLJUqPkf+jV2hii/pymS84xzgPOwmMbxfA0I3PzdDKL0+Oqq5OLvvjLYra
VJ0gwT5ybz1C+ZcDCJM5uf0j+Be21iVJRh5/mqoSXpbQPf9834wQB0xp69GuimhEURx4V94Idbmv
6/geHSXuPLvwuIF4EMW4l1piPQyRoVcGZvFEFm4A0H/ZxYILByW2m6lfapisGnEpwXwuCPA8CTJZ
WgN868bkjrjG4Xy/P/ONCSqcpQ4FzJQ4BCPteNhPn9LyMwcQYa7N/eG4IUAhRj34mkFt2qIY8iPw
1KA+A+bAFi20H/5d/5CXpuf+9LSTlCjd2Np+3zR2pqBsSS/YwvChy8OpWY3SQDgRDuuNzHRtjqY5
8v9OYnVHeonH5OKZLGaZY1WtCaq7aRemE/tCwKICG0COcHPM4ALhJR31qH+OyLBUSST8by715WM6
jsl97Lt/EsJMzCzxZ8J+MxpFjSpsDIfGx+LYZS5xKJ5Da6KPsXOuU28IBvQ/tZ9pgk9RIfp+Wk7/
mNH0QawvOcnMkIq4ycHLCdPpBBKGYHeHK8/Mi+qMIxG/jHvtfTJU/5jZMl4fwYGr4g9Kn7vbORGU
qYdUvsj4W4V6ikRpHukClTNP9WIIfZXfLFPCkBKm2/F1actMFXCw+j5zP3stwCGiVixNX+qp0VbV
b5M9osrIyWfT5IkF1FDc8UYndrGlHDhKlz9gZV61BQ6RDdIx8uBHf0RglLEru3mCA/htLc8ZX1qN
knQQyKjxbtWV+VyezmBaHE3HXCnEktl8XB1hsMxyQw7FvJLy2dg8E4iyPXdntPR14vfyi6gppp9Q
33ah7lSAocB9ulr2YqhrKZshxDmlice8CncWXoi0RQhF3kOJlOqaQHzaALhLyyf57hfmZahU2Axf
DKV/Cucn6baAytJINR2hNZrluWfwtOI0H101lKY/T22QA9X7yw3kMAB+++5McTVUzT/krKJbk5Xy
FHPERpqwuIBd3HfmSodFXYkp3TEXkD7m4Ght7QBmPy7OYSBevwen6SPSylJpK1Qx+Xd3Bfu9mE/Q
rU1cJqwU9wEU4NGtiKC/XiWDPAfp6DIFsA7CqE3fooPbGCRl7J/X0kZQVL08TgW5AVpCzmhmtuUh
GFpkFNxol6RV45hlnMHrlC/zxQqzQSOhSJI5akfXA789LThEqfXWD6sL87dGH9IRpJPq3AsGohFz
XjMfcxVl60S3vXg0V2IfpphR6G+aOQphhApDgGa8JxGZ4Hbr2XODmAmIYRx3ytqPl7Im141dOqKI
sZ7+Ui2ROWRxlgXx7lMM/3MhoH0ttsZYg04qcE8Qa+QulwcX1QhjWjrz4qETbkQKnAaaOTtqYMLp
WzKxIN6KibtVa4r1yMgH5kq/WTz03e1kw0iWtbrZOlQ/OeO1wUZZHEI8K42FGUaL0CKxMVwNADIQ
M7mvJtBTo66f8CffPdFNXCfbPa5KHJvgkRvWy0CP0nv3IJoGk22tbCWOg/2GWCj29dIrIPkE2MPW
HizusP7paMKQjI+LTtjfcRUSsFjCZ2vKf0sbjKDwQ6d+91nrTVSQz6u7gpXmH5fLEICYC1rw09tw
P9OURMFnrzVp/s/s/NHiUjzcbhXMINivCp0piZv/X9sb7oSYwE1jdY/Y9Fa8Y/ajXa0cKaa2OZlw
u1/N4r7+1V09e8LF32d/Shv64rwcm3zZvS/aq4DjwuX7PZbmqLGuGEW4i1Y28LgP7hGHxTjxkhx0
G+NfDmenYnpAnxcQXMWzz4Rk/lfc8ZwBw/zdtjxFsmJ9C1TfU9asq+e5A2juwVWPgi8gGm2MyYUF
fOX1lCQFvWMFhJiDZRxHW10hSjUVhwmq0kCmP4yOf2p0X/kMDLoRD2cUIKs7D8S3/u8dPRdwRTYo
fxvF48YKAz1LB0IhX+JpWtaSaeiughllLYVsggxGjXdW6Hpr2cPFu1sqdknzjX5j4L6cJ10gEmdm
Sm6JtZd+4/41oNpwXqT+aYbcb/F+5N4RDyB25P4unHF9OAKkUzKRpsorgEuJ1dGwZVodyixxNqNR
MAC6Pod/pVHMRJlW2q8q1Fbp6ZG/cX7hd0gXPVSyEiFt2taYtG3dOR1XfxON30oeGWwLQE7BdsjR
Soqp89xDgc5HCgrafoT7UovloOBPHj9l9mr/WKEJdtAgRKEwqJw44tacC+fQr9oL2vHEKiVO1Gvh
2QoZ/529gpulLZKFDHRwInNCI7s5ZlyttVOXnkZpRellpgm9FAo3yFuJwvkp5x0BXnhR5ze11K7C
udKI95P7Wz43WtjSRYpWyOomTUHwzEzU/jkyzovzj1eOI2//WGsBxWO00gwhMCUp1ECsklL6A5J1
iH8yYoFPOV7nJGC108wqgt9xkDvl+FRQeBeMwWflV+wItrLAg+KUsISRVLlKEjhK7XQqbItPHtuK
dJxi1t/w9qdBBkUeABdEjOVBINNQJK3dBfAE00eRKoT56caJIgtu3oIFtSsqFzhfrfOyP1VIxk1N
ghrHKX0Rb5olTSxT+Nf6QbrDdBeomqaWCxiqT9KTW73Chu/FP21jm6U8llILNtCqAZZl08I2Vdhg
tuFGv7bHT/H9wy8EVegFtS2oKit7IXl/fipMO8add895i1uq0Bygr1TaRr918zaSXBEjPw8enVmr
TPZWDsxrjfiTUNXcGQapG23Alz/0kfYKdjnuROozEA8dDrPlZxlJl2bWb5WXM6acT9OTOgIU2aAf
zXBOwERVQG2nGeT0i20MawIT6oAV4tAEZ5mpJgQxhCFYsS8qDG3vJezMSPCofs1TC02fpIh4Kgzv
yjL1AB00hNZ+TjQr6aTjVgjrLwVFLPcTVHAzXM3iLwGX1A0xH/o6/7LL7KCT0qtaDPrtZvHzExQf
ZUlT12fbiwmmGzFwHs7xyOI01oAlbmDgFUKF5vsv2g1s+ePr+QayiB7iMMOdrGMfatzo6xmn3i+3
tOmG+9IH+Aa08z3hcGAEl0+R/7fjmtYdylpLpv77h2Ur0r7nv9eOjrMRa//HxCENzBTFXPEuL5GU
NYaCHZUjWM8rOXWqbUIZAB6Bn9RCUH5DUzwYt3i/GmkM1YBl31tGuNpAkmiCM6Cs39UAphf0R6sl
W4+1wc5SKKyTnO7kEgq6AJKamN3nFries5tIGa2CjvRu5ATaUqiWJd4YkIfWw3z2JJW+iqyWnLbg
zuIKpODT3F9V1xwPbMG6jDPloyo1Yhc42QWGJ1mFj6MZTHbAzt+hCdk545CrFzMMXYa9iI9y4daq
7pvMdas8TaWFpPVPtAGgXKRRQHc9NZuS6t7rIZfHPOL2t5sVGdKjdgAGgKjkvBR78ZUosRcguFkQ
f89rQP22ynsWRzvB+RezcQLN3ZDRaxw0duAUnV5uVPrES4RlvtuHmIT14BCZ61MES1KeSGsveLga
KRqoFwX0PoHfEUzsZGjn26+Ed7RPGvF9X1B+vWqR9dLrsEbRC4asXrJLpllqu52POyNDPWQ8VQ0w
tRw+3LGznajR60AhW92pcnF3SpjDIHfq4b+czf77DPzXx0vy/vumN7vLI83W3e0pgQdddf+w4iMo
JOd18AEthsytB4ZODlS2T0ypoDZBC8NqxokmYsaetCJdBg8gg5QK2BhQ0oxD8sYGUUmFblWmeRts
q4BAUg6xutNweYKIJJcKyv8I9elziIY+T8QQTrdQG9PIfS1CaHG2Q8O1y2eDoR7LBu4Q8UPuButT
KXO99ozMHT4geq3wTwltG52+uTgfpMFBEubovxci9v2WTrr/vxn86bd3wo7CNsuyoqiOxKEJ06h6
BnevKEZ6QbuwrnH+rQOAo14y3y/3I+BTI7GlSKTmzS9xziH8jqEdOilJusIvT1rbU4KI2nvlFXX0
qzzytR1iAre2bvacCEoV5uF/9wTNp2w9ahHATP3ctupSwbsrHLHLrp3LEbuTV3Dvjv2/+kC54eEa
HwMYT5mPEJpHaspdGFTRSzaS0YEzJXbsnhTPmrIIOr7NCUc0WO+FEvu2OQQCZv8TdWavMHucakkH
qBZ6LPPUlFWxpYSXJVUfMrd1R9yX3alhUjoZGP0ptVqfwCs58KOXGHw1jdd6m6MFVrEI6tG2JGUk
l3YZ5xetB2LPb6bZERiQtMXelkZW6cLaMwm2yrFdPZytvjVMWHItymUyizWOCn4fU/QkwH/9/xhE
Kob2qPJbprqHNFsKme8wWmfZ6MJ6akztkNmNZ5qI3WZmhQRF+EDTT0QXFoYaPFAyqSUmA2ZkC5wB
2TKY5X9UP7iHQeaXDYHzKuePqlTSKIR7sXzIVuebOlmuyQIN9XEdsrHS8D+gf9O0aErRdlELbjV4
dWaJNiAIcUPAhvw/nJFhZiq86PMiUzvJ68Ve6pGBAsopGlTYrlZ63CLyPklXxTxYolP4gOoy25Tg
bKjfeYQ4iEOt6gg9JneO3Delxag7loRkrGyb/1pWaCgbhHiVu0cvPCGxF2jma1h0+ZVY8wGVjwJ7
UVtjUDhu7CdsS9Bd0UeBlyUjNNFCsK8NQW+I0vj/kPPIbMqH4CfFfz1Th91geckNrnoL6Ob+iviZ
hfxRkDTTLCapUrSZfHBS28AoWvGy5wLVb5e5z9JqBNM0g/uUlFTIT5qSMqvS10oUPVDG+zmIK4PQ
YE9CDv3YYNLj6kOmnf8i7kaT2IER1dOCOhQRv7UajCfAxKUxc9CUMCILRm8oSGKF3fldFqbQ27Zk
bnj0LUn1d9/dG4/3rIaY6PJiemCCeIHcePSA1JTlkwLJtBmgda8aPuq+uVPHD13b7gJ160dfbELK
CHb8N3ULtgpU+9HNNUqAscAqwh/q6/d8s9HDDl/SNaqnleDq4I9iJGoCfgRebMw3rfPFT3Jq7TGj
8YXWvDsaPx5L4DFGvTIwu4X9R2H31TUVDHx1acImSwBwUV3XUnyphLfwR9nR9GgxG3vqjYKBgq9K
vXpzYoV43zuAU6qAiaJfX/3UHBPeWbADT6rOf6cYvE6omc2u72GQj91G5VFQJxwpzcmtnlTfpVSa
zTng2wfkvoohRfvZzhGdPaYgT2sgmiyrUspNFzeRAqPnNlEGxl93gAY6T9hdGklY+l1TJYF2RMip
8FZSdqm2QHWhrf3TmbV/rIfyo+k3BfwNpEzzKV5KUaC4ECElkLIXmnr6fjcfUkYvttSjzZyFxrRD
guXfk30tiz2jVnLPv/nUR6DZQ2nsVGFTTxO9wSdcX7pACe3hmlPG1ZMZ/pX+9RK1G6+uYLuMnA2P
kIkziw+OXpRxuzoL0lLu2V77fiE1cLxbWs9PAfWfgtjKv0H47yubPVm4LWFRKvP1ii9vPVKP38d5
MPUA3aIGZUu6XMWgs3Q36vNuf5xOm6Jj9DuPvfuoB2y+auxeIXqnkSULWYXs5j6S6unTJX3XO4dC
fsxyObVI/Ju0GN1TYZ6ama/z8BBdss6z6cUzB+xCEOgaifdMGf29qnZv7QyNDrB0kjJEl8TAeaeT
YZd6D70f2ppYj/UsgoE64RmaOVVPCTRAZ/DCZLwVjXHb9mM+odJHk80nHHZqNU1mxF7mjUEsYr0E
yqVwrFF3YDzeDg0huLVrWlFFlUaiSpapQxCisEjCAZb1uSEu1R3N3SCiKJrNm3YBaE2OPjpaZk4i
kJAGi/6DXnJTjHNcAXIeCiNtTC+0eDL5EFZEid3CZi2F7ZdIOMTDE89Uc1HcuRy8IqZSKSmTN6Lz
FWZfbBac8J9mxO/BvZGUkFW1Pm1kZD5KpTUhcYkSPVKugZt0WIF3Q0cpHtOClV7yPbA/Dt/B0OiS
0lLT7qkK26ParwZfEESYj0ObjnT2KN2HxaBun+0DKEZ5R3cdNA1sBbTHPyiVQScNSOGQ4ITQZBWZ
UHFjkbxxSmnZwfRGQPLOhl7qWBJ5uXdcivfupsCUuKjuKSlVVojLyrvcrw6///Hc07/V/zHuY1OF
MFk4jk+IyocHQvP0Zy8oV+8IXB28vNnKUMXyM3LJ5ZrldtK77ORG+m+Z9/qRnhN2q6/eBBsp3xx/
XUmCRtIx5jcGfmuXxq6l9nHkFHzVu7EYQvbCkQtwS37gHa1+IDtWmFzmdHnJ65d0uwxhuI0R4lGU
CfjuAT1otrtwJE3INn6wbY5kNh//uXM+wn0tDgETvnz6NbBfi6vAClnsZTuq82QiZY8Ii8NckJ//
sruqn5U0Ty8kDv1Ge50SKe3WFKturBAW4nNV7ogQnMOT/Gzf56+BHpvoFW1gXNLWbubtwPw7/CIF
Wfcp2xExkJ9nYK/6sQT9gvPcL0KcmURs9UXGNN/2yhstlY3VlijsHuANExM3EO9yvFJcKwtinAVO
pXn3vIgLTGlbo1r4Mm/hnM+BZmFg2kQWK1BE+K56CxS956G0OK/J/31cKHf5Mg853nDYnMJQcl5a
s8JwA4c8hsAvIKFkAYZ0xMurD6dUl4KTFrVf4iyg0tTtiqOk4L7gqj1SL+D+ZhX2T1PYzj1yKOx1
3EuMGFezajZJuY2QXuOqk7sEux2qQF+K5y4MNwZNz5nZK0fyrSXGRI0JTpxQVj39GZV7kLMKIL7w
Ygwj5kzu5ZGd+BM6H00J04hE0iXdcafSLgWC0o7pddJsuY1NEnw2fo2dkhbFYBTqKnCxnAMXp4TI
dhOh4XrxkDFTf0LuHb3xiJ/YteXdUOeqGEfnHQh++UkZbr/BZnhq5+9m0ycLNjh6xSMlazM5Sgtb
FOTwC1MK5nuwbgdTg//k6/kNr/SqKBNwyb6rXEkaZ5Y2DSBaj7mGBdh+CyuJuN/ZKsfbEDv0XTkW
qoxtqZ/X58cDMDof0S6Fu7V1gk5fo6vM42G9iAX+b/tChmQ52o5Iqydalpw1GlLZVgAlvCu6R2LE
qyGf0Rc/TAlt4ek2diNI41rk6Csn/1aLm8K++CyX2TmN+yvz0ox1amB3KMyCnldxvjBRMKX7oMn3
yaWt0PgV0F90xFnxTlkrgTm+AO0rDW1Rnzu/u4Q3dmUqCXaxpsG+yifgMBYuUtRGZmE8vUGn5f0w
NfDDoLi537rL4v1fhpxW3+jVQg4bcVjApdupV/+lq2VyqySCHFpcAbKck4RROcpMLFRJMdNNhPCL
q6QwZy2pZIJ3kFFcVpEyE0bPJKRHCK7yXEZMfjTDuXwCsGmMYvaegNFEs6RaK09i7RXO+sh77bRA
c9qSoofQjKxVLMaFgLtIQcDQXa3a+nQlBwspAHsqSzBmNdY7xBh2jNBB1ThTbWW/WrzHKdrnSJYE
I+9N8C3WZPL4ix9raxyb4II9HOFf33Z9L3nGiMixShGLTZkWIccIZKh/N7lfmrYIMIJLiHuMcr3n
N7OR3RxTokTAqZPQzattwTN7Y7dEUm8L9eSub7chWiLONiTAc5PQV5uwsfY9uyczKIdBfhbQEZCT
fn4GYJPpH1VgEPSWm6m/c3yJpkk+Ff0i+S+6nYRS5Qt6c/gpIYBK/+FCNBtY5aifmRYBJKajtpkW
9n+zp4FGk04Ub9Ky533figF1SQgaGkxnRrw4R3xyhMW98IOB1BILEwGZ4THKE7k3Nr4VjnTEcziq
l1Psk6G5ClpxnersMTrOV8GeKb/mADjgbtph1hW9BXTiAhTgociJmZ4NiyI49IYveoP63jwsju61
Ss/gLJqHqe+cS6cza5LkMdNRoCecyZx83k9fYSkXM+Z5sHfX1BA5mHxvKkxSjiAdCuag2jyXRN8Z
/+rHPaglB3aLUPQjW+uhcy2psyrnJZkG1V9Md2E/5k1JVQNstRJ60HkYD58kesN0uHGbHHbqVd3U
FKfOcRkWi7kpMRhtcZhqhovvTa5KyLnRUzxzjR+x2MmNKPRnyFIz8MHmI4tHgtMNVLSsgY2jPyGY
FvSAm9yW/HkVi2FB9jfYKdVnsKk+HD/GTtIQNFJ+enmGrw5ahxdq5hIaBe1CF684zjlQNuSVnQve
oPLY/2gvSxG3/aYZO+QmFsqm7DDFkLcjv56bcKZ1+Dm9Y7LVmlsm7FVvzvSHfDd4+V6PWHnM7r5h
N7CWEvXk8KpBi3bn1Yjz6lHHJRyDMaePVQJ1zguxZeEgOBMIdDRMn9ELZ3f/U6xE8cUUC/xd8qoY
u2Htx4F6Xf0lJd5SZGg9k3gja1ubxtPRdD+JAQF21KsP78mkSiZZWWGwY7XCFNxkb63Clc2zsHT0
N/EpBzsxbCJAbuHNdBHFkuWjt4Kl7rbhYMoV6YA60fdvSgZZ8r1idRyTiY0TLmGiXTI+FFqPXm1V
Lx6f2Hbe5SIQ2Z02Sf349ENqjLx5GI3vPt9NAeTqVQlh/jPqcRtGCXBUojG8Pvg7uP/rr5sqayOz
EiQIUO04k1ornmcPFgUoqyxsGXFwmS8sjdiXQ6WI7Djf2OEJF8O+EQXu0jhDAT8hm667oJjnINXD
WhxzUO+Knj3mK4IwG3aPZxiZvMPOqXid3jwmtIRDbpaDuvk8ibrKYGBmWGagDMIfSA8Iarhugd87
NFI7EluNRxY/gdpHLKpd1QyApu6Puxpo2yDEcoB442huZ3Ab6UMHXFtzLm4wD0uj/5Tcn7Rx/aZU
EL5HHBYgcjfqmw+Byn+N2Y5wBWT0cmaYMdwTpid9wAcLKwydxalJBdvhtZYcHKzhjB+HvQemoMEQ
dE2dB9wRzTUgEUCH8TKDYUHYwZEimg/UbuymjsbOaIOK39iLh7v9D+p/kGrwLyg+BvOaJKWOODrR
oxMurssi5OF70sZQfpUc7o/BMhLrcGuIAFXM69VYYyYESF/QJ/4d9dfvaB0GpKy/VWlx3q2P6aDq
p2LWL9XYFg6FNe5sCH3tMYXXE2UM0h/DuytqubgViZwdCmy0NIJQXFos3aYhnRwCkpUfDK+rflKg
qZP0gUwT3gyt0PSaaTgzBB6iaPYi4R1Wj6fTXTotb283O9SBtbRUT1JCNk2DC0YJG0/7CGLMDcn4
U+qaIkP1IgGiNbtY+IuZZIqle1HSVvn9/VuiEH+UgssJi2e7K793u0yss1EqbhJrobqFh4IJr1N7
OQaNuRfZwJYJkCaJPxeoDlSQxeCgZdldXXUwIwKW6gnWgJz/YBda692A9hjY/qvwaKXYfkuGnw19
NtjkqFTIJw3vn/nhmLe68XvlRTJAbZ4i+eydt7Z5sMkDrWkjPfwmaQf3QFyBUYflVOpW9jNyGhH0
DW6uEmmp5iIvCKkSx8O7iuGdGJTyx/XdV526uQbX8B6JBiGcPHCFiS1TCYT3DH8FajzG349ZWri9
na3iHdx8NrQy79G5W0vH0hfucZD5Twvs/tMn3bNsAg5ZgjZcPIBH9eFB73z5lOBIxuxRV3CCdjQj
zoRzAPE1V/47D16XV/zzezyqdwlujqMtdt1KXArnpgKlZmyKd8Xq4+UNT+WisKJuPR0yUut6NvPa
maCzaBtLRLxNJoOY+zbB7dsVlifGbp2kM95QqrbGF5bO8NFDwLcGDeIyDwBV1ZoKuJwmbbyvr/lo
yJMTW/p2BnxyM3QCrygx07hr0ClHqwfI+U0E1i3u1z4JT0YX9d6t4RusUxiWMIURkij12wVrVC58
vJYy3kQtwRRDK0Q9J3v1QhMeNIoRyRTuQEB6/1tmgAA8l8VH8br02YobdsMJlJiMwykbpy+lZhve
Z6zUVpQbK5MVIKVcmFXYQxYbfXVPgq7AYdH5NU9llJjGW0Po27EGiTGthUYhJwT3bzgwJ0rKIZ5t
zJZWpvjOXcztY+/g6DwGU+VTKSsB60wNjzC2IMh87jzlWqD39Gyo/sYiK8QMTWuHemXXVmXes5qV
S7TAfbr66SB/rSKQVmmsHM0/WViVwbGnVahj/7diyl4FSNF9AQVSCUQUjeUBMik3Z6xzlA9QE3zs
Ilhry37XVVO12sdDvVKIUtAOeo4tf3vFrxnFGjHueirBHI8idZtwDn58GtrvEz+O2Oo9lqRlfLZJ
uF65fNtr5FJZO/K6hL1rELTy/vwdr4ZKOKwWk+8qZ8KcZbz/KlOP4xAd8k5WuhXEvFzYNRziW2J7
6HeVGdY/ml/eNq94A8wOSQSbGoaX6plw00JOI1ClzOmTSYx9yi+T1MLjYoURdlxJbF9wfwFABNGf
CJOPE6LWZVyGSkXzfRtpBXBv2Rqerrrd8e9poOBYBoItJz1xMG2XaG1By/GW8qRLRxnvHaMTeDB7
Hxn4JjAX670g46gURUMRIqNuKSo/fiWIu8k6R+dkUkMYaW6exPLQg7xbR2a9Zp6Bd8Am5PO9ToYT
MOpWniWvEWqer3Hy+cvvBIQ2y0EIEP52N6JamSoW7QnobOeaR79UtNlOdsw5dTP+nei6J4vZsp3b
LCsDi5j5L6wRUdL0Tzs9RAs81zXJMA17pBVjkG9Jmd5V0sCMo0jl/1HAKKcRBtza9NUkt2r+cGsL
SoLAKnRX//0G5KCEb93IzNy0HIj5p5ZqFVs2OAMh5JQjNNZKMVfz2grHT1BMsYnlauxiE+I5+7SL
6lotITZGkMfRMvx+YEbtq0nGh+EzZ7lbMCMl4IB97Z8wBgHvWvqGhPAQOW+tefKWQ4qqBHf9vyGs
JBEf95k5TnFtFefzrtXHEcyvY2KOPFrnv7umLyRZEF54uCpIoU/XrPQc0RX0VAqYvT0fcpcg3/9f
fCZXBi2G1lQcIGqZO3vFaZGf/dOCXRfpr+WGjUPyN8ytgehOUJGYN8hdP6o2bs4Yd9YmN7TmKJQs
N35zUOJxFLZYKnDJYjC931SqbQnSgexRNgfdqyXMhX5XVWejyTYgQAtqp7jsz8TiFOGzJcxSQCq+
ULyPERu/s7EDQLIj7cyElAXfEPE2sqEDGuh/mVwblyZXVc8FU/UQghAqZgWtNbY2NGlcnQ2PSz/O
G5yrLwE+uBHUTTxtVwEpoX6iiNsD1t/irNfYLcS9k3XgSdFYUoOB1+eXgBWcIzYZ76tLqjc75OTC
EbwPSF0kNkt3UPwyJGLqkYWh874P/4JSTHbacXgcVvvubIBiNXr73l6FRnPiqpvXUFXKfXEHcS2m
IoXMDLYsT0LQJrgiWauI16S2/g7VIyj6/QVJa2A1kl88ugqWKfHFOe4ZXJRHRS9ur9ucPFrKNg/t
0iVbth/mJgK1F1Uaaf27pShUx11d3J7x23fzjhHnPNjmz52zFhgmqhttEVuHNc8ZPhTScKCFU5DC
pAWKoUFnG5Se5AbONddhXnS2onPPRioMA7Aod6X7jlSm4aX8aS3YYg7y/D5imcyMX7rlnhQLwShk
v784RpIZk2m5d+0CYrPd4k8f1/T0BtAUjyRjYcB5/XNTu/hJPD2xwAUc8DaBmsfsvp+LyW7b8pIl
OXcvfd/gqLbPWBxtk77KFNJcmgQ1paf0kNjNmIqflJrRn+hzC7iifz8ZbK6OzT8P8RQyWEdWWnhg
Yr7/E+ZB4tytidfu73Ts256ga2JAF2KGx/h33tvE2UmlnWBCZbHn5acJvsGHrA3AgjQ8S2iyOmlT
+FAAUPsayEqzf//MhJYn2w5Qht2Sb+6r01pPNTd1grT3ft0C4rlyjQzPkoZiP+5x7POHggyMIXmo
Yt8Pa9Z4Xhq7vJ2IWq9vEZBs+ZylOPQkOmBLG3/6WCoX83xaQueGaZvCIrYBPqJRUvq6SjaFfIyA
NPtQSJitqYmJg6/eCDW+8Grf69iKBxojJtqXuVbkIUc4gFq5DJOBXZUHpXY7f5tvqW25rrYE98Ec
keZiwp37f0tx9o21941TMBDGaJFTdQ6m0TxXWKt2n5/+Y77WhGWQM3M27/DNQN5qrX8N/6TrH9Io
Tfi2PKaIYLsP4N0rh1bIOIQIHVPNGiiFv56eiiLNNop3XVhLHcGQTf0pcBgPWTgUIjTTjrBMZYNE
S7g2Fza7qUv6GLl/D1jXoXawfFfttTEohObRaBMyR2fa2YWlDuXop4AAI7qeJW33YPXALX2bLdNH
ByxtnWg3GI5TsHeKtX0InIM/TJ0aRsUFETOnyztKFa3bTNmVIu2IvEHLwN0DpDFHPIsajRjKMbsR
mUtC2RRyBEPud2b62E8aiMjsc8TCNgSRGJd2zXvdkzur2YpVKOrWNdYLEUMLZsgW+ixg68+v06oJ
F3stftOWxD4OMb3y6VmRpUJJgwBOxMWWUauadFrVEa7sOcKvOfSDYM6rHIwI6NLoUfWUK7+Vc1Ma
23uIRmmCGJCH60V6jWhCIrnlW6LnRFZFWlxwaaHXbExFqcepfOF9HKeJ5rpDPGvr31qrceVyEngH
HipvFzWHQH93alYNhRycFGUNwkd9nuVj/+IS+1gFcAs5zds4BeBd6Uf+nR+AirndyHObYXbf6NwE
yILFH1gy5Aas0N+LxdDRzMOsWUNTXh4rEo77EEpGuwgKRNeAs3MCrk4agMva/gbDozS0Cj7uY6o0
Vo7mo5bgGiB/LwpbhVv/RFQspF8fbvgPfO58wmn5VOPaqlRf89uR2FUQIVKJXuFDlyG2/cm+Na1K
F6NEEF1gFt4e7xMviAA6VY/EuE5SHQAxpeYozljFC2NdjKJyES18l8QPeR91NV0GXHo7lm3kWaqC
bLVfIxdorP9xogbJoOaBKOYwCrqFU5sfzIjs+kqms3orbPDwatzkrXUWFVNH+EDMrAIB6jcybl1k
mbz1Y/mvnm/7klOEw+UibKiiQ8ifscCa71hCK9x54Yboi5QNNUfk8+1QrUSODrD+4JRaoRwum6qr
VhyM9WdSZ0QKUYurlrGnj/DoDqqsudFzS7tMQXj/B4BKIMTRELgPjHrwViEXYwYWZaql3FZd+imW
nbSc0I4m9XGUvdb/JMsORVv75QGqc+oTYdKQaqeswvgdl1UgCfu4xhURVmmPHVQziRsYfRF043tQ
DMRml+YoUeHG+bJaMWpMd8cXpxvvjNiDDttDuym7LgvqacKGYvo04HRDhp4Fq6/1GW1xLFoFI0L+
kXleDvot6kkXSnlEvzDZdHpk8UIDnq4SHzOrygq334C3ODALUqbyLwE6XcR28SG9fV52HdbTCn9w
QktRpG3t7A7lCA2WwDKq78WpctDHSVL/lsw3GQf7jQGTMeuNv0tcClySAQ/HuHBIl6p1smRt+akT
mC6COp9k4WY3awWUozrIH0vkYWt/2PTWlJm2aD0TGHuZoBAk+BDxyAoGw2BX3mxKgmeTYWyYzOL6
4LHtKpUKi7BHbAsYIVXvhML0nbUgPDqEO1MA5j6OHy0pG83l9V9nHd1tsnPOIOjLdJaD5noKnw1X
SptgGg4B2Vkd15xoe3nGEcPTUS+kBXp5XoaOFAIwQyVG17ENrbe1b0fZW1lMpc+aHiv8gFzcHQrX
Dsln9nmdp7yX+h0uxE++pS6vPRbBuyXPH1Ronybw0kjQ4RC/aohyqTxI4PuY21WUhCgz1y0BTOTl
qsZhGgKBVeA4lMRu+kEeg9YOdjsFkqUy1Y2FPEx0rkwxiVecpCd1zSkQQvEaU1EcDHAyjcq8hE8q
o5bE7AIYoW6qzd5ReMMTs1MtfEHhtK5zQBVDDZlV2TRRAAd45xYjOrJpO4AqgRiHk8IUccaZf03w
4Dt0lXS7DHdpMI1W0VnBoBXAn4lLxr77w94ywdjl4x5weq+AZNkQrbTBCQre9ZKP7vrk3Vxn3LTq
ICiO6O0fl+8eMDbrp4yXVqmUAXm+FogzpVocz5FhW3L1sU1Jy53lgban6pXKDwj1LyRWUBxm53ZJ
zk4JYagzthQ17Je30FhMBANgrBpp2/0tQRuCPHJi8JODcN/Mh/TrzjoJsWaY9cNgF+XshC0MGZn+
nDhxTgaNO/CkmLt017g/DIPfHZ+QB/PKcLPbk2YuehTSiFXVMh9WutUDRPqSuAumR/nTD6KLAbgj
YnXdt14a8x5Lz6FR7xUpdF11j8kAd9Om1GXGcB03vN7kpwoBZgDn/O3sUFkQariQazntJDyOaRmG
youTICFzACzVC3MvE7tNKJLmLrkUpJcWSVRi662zElFC6gSDh67cXrgOVGPiVT3p98uPxhZbU2LO
0VEqcx9ABaxwdYxKANoH88/RaeusOkgDJFXYzBTpcMHVWHKZ6UAYbC5508CSO55Gt+WnWIiOHByP
3qYs3XzvZBTHjvB61+yrylvXYCWqS67WVvPzf7Y3VBFj/PbmnE+KUjOqcnTpK5n6bFO2dJXuQoG6
q2z2qfYpoodlgHPk7FSk8U5jkV4pjffJAkI7xmHqmYerzTQO5/97vUS0fstyijcl7nQnOkaUVwec
ZwmCozBPVZ9FCEOm7LxO0GhaSYBodOE8cQKJ+lY/ns1+ABBZ9d2G6SPthmemPy20FYi75iFh0oJ1
JtbwyXMnLmj/3cglVqtOKYX+gQdYmKBHuRP5SR1xlq/I7qhhfsayYwzhQo1dXTV1vst/fe5eHXmH
ByiY4A+KSmX0WLd16EFfY0cInf38TvyFgXdZPqUNH8Rdp3mesov5x1ummSSoIOj7HM7W4rkuQJSN
7JO57+mxGR/AJR7BjPkFJC9Ho2hU47iKpCk7AANDqbvUKO51Jjo9DLQZRYWJD0mUQtSnKmgF8s8V
tr5oQEFVfZu/bBWSTTSJeXwDDK08zKv+GD+QStTusTfiWIiF5utXgJE6mkN2WspxejGwpcZigpZz
vzdltC+1OfeUqZdIbXymmd60dC9hG0vCG0uS5IIGjLjyJcA0bzdUxWEUigJ6OpHNsOVx3TM5Ob1m
YrGyOJWzXG+GtQ81F/QBCdQQlHJfeC3AlyvVsNdExKrUWAxhp0woirAHFlU3GNo87aK67FcYTMMd
ls32JXALGo5/8xI0YXMHZ6h8LGQE6a5WUwXqNatoRyDKI2uTjJ907ZMIRuKj5dhWZ3Q9XTMroEJj
M6+hLV3GGZaXThsAZO+B9+VwVmXl4kO0XA/tmL9rrCmzahTmcX8BAe/Ra8Q5IOIduLVcfcOmjpyy
hjuJ2LaUjhLmRjg/vQQVR8cIAixJKQj9DF6zumgIOmOBW8iXnO4LpdR9FgXkbILq6KH+DxSo+hfK
zQtQblUclv9yVdAhj9htatjNKjyYxmJc0Kn+xFczuuYuVuIT7fW3tT3uP/KwmLmxFMShhxOzmumf
0LaSJ81EmLQR/K4ojog20Q63CfV830c0g55wJosM8e15ZBAnNiWqiwGUfTuqE2G2VNbVQtaHfCN/
oj+xkdl6ut+Fyl5KekL2hdOzljIEnBraKhd9Ief0isgeKLYuxuJKnHsBTbGm1YSKil0KkENzgXf+
j0vzd2xqOaM1hONDKC/x5ic8kidN9krF5SDpHoSEaMU9azNOxwxgIKBFt+Kf9oG/h/gi7a09eKtn
j1V6CqWVUGRxE9Qd5pcdc6u+KCAP7jgOhCXW6Ppg2MRF+ZasAAKln3BFWvBzdQZmXnbLjo9lpd4x
SQTmF8DpApuh7aOK1fWiMapY2Mlsyyn4ksqivvYP2YnjR2v+IZGmr8f2di7EN6sBZdQXrL+5MNR4
VVQ6iC22zUSg4r7nL9DRlr9L36PhCkjNDe2CSdipiKHpQrsJIkuNigF836e5e62NTO/G6yQ1xZ/D
sduxluRBnpwyofSN2en/EX+XXcCaLFiqbPRw5ruBWQ3hyOKEjaQtEqEuJISR2DsD1RWqZZUL40UE
982IVcyY62HjKf046NW7z6cJpWYk78seWnaXksQ3zuiscIaxSHoWzOpRSVhKYwdp9A2ljI2BJDei
jQWw9SBzj+rynA69loNrGHuEmlCtA2ULtgeUdMO4kJEGGqBZxqjXXDAFFjKgN+ygjipnL8WoWY0r
A7V2bB8a56dXZ7aORt/+jwGsePIoaDDaE0dKed8fE2vKD3EuN75sRtZk22GNAm8dKniP64ZGBzny
/p++eyEZwzblaywR6Qq2+8rwAqyN4xZAvupE+v58M+NW/G5lA9V6spTBGNN7I/KmtytJ1mGh18ej
vtjBYeZ1YFgPsfBvAPvdYZyQRWY+BHwwRuRhkom/cV+3431UezhgCsHn1lUTjAIX2LCKRX7dm8cI
2EgEy1evRoWW5hYBxospjtO6cKd23HGHpTp1pY7CCyInq4K4Daxs1Md2eQyYtwesedpFBwG++p6a
dU024ujDJcyW+MhiuKT9LcZdAULvS06HE0ZmQBozqGhHi0sH2xzWdy6RGnsPNjBJAPr+TvBHYb4P
/G0SVeVPYE1inIJMwaEawWo9LuYgoLG0HMJyGfkTN5g3Cg19qR+2MjgaisMUXgiBjVnSMLhLr8NH
2Q70BiU3j3cujIFdq/0B+uTVSYuDzhmZG/zbnZ/8YY+Sf2GrBBPyFLtbZ8Z7sSNTxk7QT620t5q4
JGklu6aPGuqrADWpx7CBQunXyg7bIjPPgEiUhfp8ltyXFA20hBfXP248OnxcFwwUCjgaxMO+3j10
CMfv/2VmZMFNDTF2/j1NRTmY6c6gS9rktftqxhB/Za+RBE6EdpWmCr4+Vm3OS8C2VhLOVrfZJrBF
JX4AB4oaUqM9C1fd9//VzXmOU2hDKVrlQm1qgjelmebJkFMeLzi68G8M3+rt3zvKBpt2dPSAZjJU
c/7KWIXt1vvTF19uW2CeNg+29eehx1+jQd0xFOZ5VWi36q137TPCKL7nfcME/M3qNFxtdpzYTsWV
pj+/3PL1d0tzn227iLM+WnMB+/asSsxzzMzQPe0XUdRezwO0TW4hpF+JQcAQfvhReksiX2CkiYB/
FYK+Tlu5mxucrYrbW6Fkg/9/rPW/wDik5oh1H9y0rrJOUEBvBjyqwkMja3+3yYcgg/HP91RTWOOH
PR11HSYc6Af/pFZtPLp/OQLcveP7WEeDu6YQ6QFPv1E9dGyDMf7kBZqzW3yIWoSupZl9oeJpVOcB
MsBigEGE8p4xWbD1kmMlJMud/+inbxR3lurL+aOHdIa/Nb1eVeEFwfAd3eGTzZVrz2sA4eR/bJZU
KzzY37LTW2NPsNu+vaJtt/q2zbWvuzMrOcygOutUEQEzaD+HKLsuzjuArOo/YU9BE7gAfEGJk5s2
F607+uOlmxsWWqKtxquTDvgiWVzQSF1PT+YkO1Q2wdur+5wTFVW0IqhizM5Jss57CsKJ8B/vpMdC
es5iVG41Fb81NQYXdJRAj7WVCCkt8MNrBxGxhg/FDkuYTkw0jHiT4yXV703At/9eZ8+7zUEPbU/M
tpRXJNUevwFfgTSfZf2d0HwhmIZ6jiMrbOwyy8dnNTxVzF1+BxHuMNO59WUK0vPOLIthBQDZ2Mqd
rPCQqTJGEEa8p4RznlhojJ0NxMW2om8DWpsektiGusZ0tElfdKFhCdfWgd0tPEFuUnQxHVyjsQ3r
eBwNj2A4yZaHThgnVs2zejD6JBqYoIKJUo8zuITIAhPpv/sPRTDlJ4dsJr5nS2QaAZlxMVfsZa6b
9vq2nsu9FoNGcqyuB7Nl9WCY3u7P2nJV86dGhq+X1cI1MFydY+zPxOMSDSm/iFPp2HlMiG6a0ovc
5o7y4QeLLWfO2e2HZfkrsnb+LAHRtdV+vdteFC28C9eKknqre0D372yRTqXx56QxNSbjQjoqCOkq
4pkfIP97d87p6GerMDlUb0eNnd4ztQYDW0yJDvBRlJmuknMwL8dWdXbaiFLE7Zz8xBSr+L/KmcXr
tZNXM5rF+4cJaR+63zXQjwl7cqWU+51tEC5FJiXUPWXmsmle/vGoQN38tyszsZa3WjDPxgVZGG/S
gwyG6T4acgLzBnZyoydmpudpGcMMZFZGN6c4S34jCT400BLcrcylbd2aSZr4PqrAhXyNQL4bIgFU
Y6sIlY9s3dRFEuHIgkRoPEzI/AoTiCfBeUlIQ5Fs4G8PQmRkbOdjhISR7ISwyox8LVQ9wSTdn8mI
8/g3WlkcpZgUYa9BMLKBgvrTmp6ez06Nu3/TKKOtRJ47jINE84Z/6MeL9QPRKy45sHDMpdx8JqQ0
hFtU/ByOPiqbl+FmWlijvel9byfFrA3TqHjRWOuF2CRoXA9ASd5ImtMW89oS7Y2eJs7Za1zfQVtM
QGxZWVWgpQCQLbAAyTFClphp8qlUfzyENKlzGxr2ic7AeOOqY4v+T/qEKYvOENgPPbekzdTcfx7+
ojlR0FwMIk7be3ZXDxyDUO7KLz9w0WE8aG4jltPywvL8+SSxSfpsqhHLmvTzUYyE6KQ7rEo4faI/
J8BGL5jlSOR2Qk8FZE7WzgdYQcwRSyDOXktT9Wl/yH0oGzssBg9qA6qN5ZWLfQgoEoAp7x879x0/
4b2V67esvtYRChyR3Veor6o50tC0ymAMXH85TvE/qFCrdR4FU4bLv8fR8pb9/RJ0leQQWvfIoUIa
hk6HoqRXbh30/Q5jrSTCtZU30geyGsmGIthbtNWo0fOakqMLKGxQHibthfXcY4KETydt5R7gneNV
HH0vvlgqVp11gY/bvCNFFMOzhuW2AVm4PSnLp2h/hXhtrGwGFdMIu7n44VYkMchLHm3g5SnqFZEr
kykOQ+HoZ1hDVv8rOLXHHVSZJIPLyGYIELQBTkPd1WXeMnR9mt6Uieo7UPVwJIh6Lwu2Y1QQ3Qgk
9nPEU4nKpGeC5CQ4XC/8t7Vx/0mtPbUlUnRNfn2Z4UHnQDd/DoMaoHsru+VOCE19A4k/cwPpC/wf
5F7LrtfLBSR1svCvkkQot8ZSYFNFZd0a9gjU2Dxh05DCoE7qqt9fL7PY/zfV3LUGlysIutO+oGFA
TA1/6Kqe2zsMvQhPVbXAeo595Wnc5AY2AMzfLlvWmLeBmT1osUXTxh3Mlyb0dk4DYEvF+rZ+akgf
5bY44fCCPIj/gtwcd9O5lNcWA+gf8Tay8Bi83NP8CfoOZ35Pq+KwIFVftQ6xdV90unsDa8a8DXNd
rtk/K4aQsaoMaMX3OApO919Eyle240vNQ6L3wWKLFYmuL7hKchPx9ZcYmtpCMVzz683/Ux+Rh59Z
ja3k0WRL7epK85kHYxEumto7PfqIHGW/w5HwXxeuDuBr6VjZiFmnOePX24H4G1Dp8U+OwDIbl1AX
jdSnwNF6qkjyLPTD317nhhrlJPun3btbyHgGjuR1bYwB3BBTvYwPOZJ6X3SFR3atl9UlX6spX9Cj
nc5nIgZerLetb3e29PQNUlKBmGX3oYtLZ75xkhmQdqhl4pHlSgtVKOAnJOKDi67FSx0OL2MnVdEc
2uwq2SPdkNEn+6DKJ4K60VmVQryahtl/6n+Q6GTbxnM3nZ82IOWGfaRKATm+FJtpseAZCA8GO+pP
z2komZWQmElKAkQ3MGNWftgvMngP9/XiHOLcgx9rHMwmML8Q2JhAcDjdYPFcFGYO2e0Mnh/18x+X
b3u8mgggsxYLyRGIaj8i8s1DSSgkhBsr9YdF+C/tEzjfpKyUzUvdg0soqiZNf9HI8YGmBkJxfUqk
f4wfo8gQkQZ3D2kbOHRKi88yDChLOFMyC7gRW3z8O3KfbLFXsuo9WicQKUMOqAlDUWRvNy8dJOBe
EqqTx4fIYvN6o7GeJgAdqYywrvhZAf3m+0+3lGUZnBR/xE0kwDtGplqKneb6DXLdCoTi+hQHW9Jh
+2ykSCkTh/Egcws2B7qciHOkQ4daVTG3d2saa7VsBD+k6Jn/Wld7ebmUxGPui9eSeg5jAkj9aGK7
GyolowdnZSeBODir6DUXNecCWAdFiXwYVCZqUwRk/iZmLrPadfe3eTjG0hBf0jDLqZtYQW2FUG/Z
Xke2FNaoYS68e2lk/S6y17i/PCyZd6qNFcKHr+PL993V+rboE+RIuj/6/Ke9b47hIjFDVds6hOpz
A+hSup/EMM7fShBKCq9V/cb2ZnhEh5PxuzF7l+63elFbxeGgDwH818m8bn7fR3by+D+xWJg7SqPB
2uGoCpn3DVrFcXh/n7n4jQdVmY07/RqC8/gEWelOMEkBlQxWkChWtvI0x01m/BIVQ2zjgA+KtJaL
3Z60dpOFNXdqickSd0yPMuzPzWE7wLTra4nOtuxkjfrMZUEO1oqoaNDpR5Ff3GjoeeBOiYlm+grb
XqNYgAFx7exeSNluZobJTXll/2l+LHoejyvmySb4nsU33tMPbfo2zS8VXj0iv8QI6hC0+nBklDaH
vFTiq/Bvdo3W5op//RmR5zjpXb0FCTjcWbfWdNJCUSPPYH45kvYUtvnWE4Gw2uoXfwjxrf8cb+5p
ALEoPpAKn3uIXVR8ViTYoqLCDJ/meHuYTRAFduJ6ODyEt++JMWZnO3442l2wWyZcoNpI7UHmYueq
0+5I5dp3Dt7ZJZ/r+RfaUo8NYDiCaDTMv12v0D1FEiaKoQOT1UHnTuzo/77h3OopMoFm4I06tNwz
ebQkJMis32Hjm5VgNddtK+CKBR4Eq96prTWZisqTFIMkmsjOBg98Xulf+bsFf+WgAy+w0y0o0LN0
zNTIe6xrCraz/N401xyAHfK/NhzbNOFunmg/Dl6UQtAeRotFCWTj8KNxJJPUnnPkcn3wCgtM3aZl
Y2Oiyz06mjKYTQzmPLXZRrqC0rugtjZGQUYF80Ly/VOC6YsccYBvzNh2XcoCGWWGbFl3t9ZJEj77
HTdIgajE8pJdORe/1liO5+9yxzy65HuepIhsmZQvEI6BbQRMhhAWcUh7KCI8+2VczQUD4ummiXE2
ghHWoV8EPQ0U4RDi2Z63zcHUrJrka4pGluQIyQY+Jwa8QyMeOOhO4XHUQEdOwIqslUNcQI3IToIP
wDnqQKYrCF24Riy2R1+vx6a4o09Whe5fQ2/4R25wT8gZAFeAh1EB988j0NMgwThkn5efsLF5+g3u
mf+cmA7GkUWEdO1Tkrkcr2lq9JBU7hjtsNZF09PHkgNRs45B+Hu40LUZ5qZ8c4z1nb8Ye9rgSokF
8IwqC4qm3/mRQ7+LhVCDSY2XhPPG0VktnYkIiGJLrPU3ogVaT+En1rNI6Y9LDoAL/GVGE7EJzhIA
5MkFzZSKaWFZqFT7apAxktsIsLdqXRBFcxQoc0M9QC2BV4PZbUjb4dACPv4JZt3l9gi6Ei9O0Gk9
Ffp5HKUaPPFN72oKSi2Jx7mX/dJNxIF95Nt7gbarRbcS4JxQKHHnrCSqJo0PksfUQINCi2UkaqLm
oXxrwk0mUV9Oj3td93p7LaQfK/Q0MfSCqbTRmz3+uEhkS2SPGKIm86cpbsCxhtKX58XyFZ6xFB//
w3d0JfLZm4uDZbSO7gUKdibwmjT+gNBjL3PQ/GqRtPT2UyLyKoPF8huiZCg7VGVgXxOqx/NG7ANx
IDQc/V+lgCShh8jTSYAQ/LhDGTenmzbjH503AbaW+FA1IUZhSiG0dxFJ4tbFVYQ8x8U4v+ufv9aO
ulzPF0YazmkW5j0kbzu6568LXf5dQnv4JV2Mt3YXTzPX83JHFpbT1VglCrUUvThGy60rLCPtROuj
3no9QFg0WncHI7QqavktcZbyGDEJ4Mc97d10yIaoZw8uCgDQO0RS3HdA5jYF8u233wq6jLGSi0vv
cgYuPCeXk9gK3W9hYRYNiavKnrYZAqGoXCxVtxixX7OnnGIAOAFC6XBBv8FRE4bV3UhGtIt+b6aV
Y8uddeLJYkaIA3gDu3M6PsjqlaNeVNW1+lyVbdZrvwhgYZB/zBEdOz0/dsNCoVSUxnp/LtKSQRO+
0HcR2JHR5rFVT8mm7BvCARWcCkZbtmUPuWWuS+jdoqsT6bRWX19OEWVY0lkbOWSiQc682BsVt5MO
d7TMiwno4yvv4I0JBE3W+1yvA1QtHBv0YwjgE7iOSpP3lyxyNljBfzdF+n9E81fdmOlwCAGHZVPU
tHDBqXZg0qvnzQujPn0a+RuM0j18/iZgiPKUerQtuGg5HXrrfwQgbT7wn9Qqhs+QL4V7rUqlgfsV
zLV5KxeWqCdUXRwej02aWqyNakLKbLH4MBblruy+oYL9kZJAjE1L2PVUhuwwvkP+hYeTtfnMXNEG
297QFcOBqn2trRHulfHf8SbeADyy6wSX4UKGYhSW3mBSMoLZf905UYYAiQ+EwjRwD5zceGqrw5o0
LB+z1S2uJhnmDDxcJb4NZwVHCRHJyiTSIH6FZXEliS7maH/SoFcSjU7cRZKCnNw7qiG0+KFZL+bf
MNacBgy0OobuXh99rUTu5+rsZ/gdIagUJUNs6gxuami6Jqtoen0JY8OkOPjaLn0db1Dz1ymEvlPx
pVm8lN05SDqXxp1GXxpSCevf812TawALvLHDCTlQfSlxMqDQ8VWrp6pVWi5yfVE1MXuISARRDVHf
U8vzvx3zdXr6lxuB5KkGUbDK1+oSOrqxRXBCLya1Ws+XQDelcQqiTuRPk3WBmzkzPAQPqQtycrWQ
H0T3M0Jjp7xW1dCRZu5Cy/fJrP3ulM7V/Bh94jzRabHthrAo0grMBQW/IZXF/mEW1Z7xBMU2oOh8
3w24WJfD3cJ5III65ivPNT+KoENhI0Wh+R1gWlQfAneMuaqRE3ky1SZp8t/q+5S9U/+gflHS7T0w
4DDj9NNtTJV/T6tqN2L7+XwgAT0nR1qBi7+jjr3bxZ0nqmZr/EpDEsr7iTocmQO62mFGHRvWhlpS
/TLYh1y8XGcyZFNSSJPjz7xpl5DLeD66/lxtY9FbAaH6bVw8R/Kq20VCaxtlqfvB2ldlBm7j6Ke7
uqg0wooSWkt7pI+P+AJUIJIP8+1G6RnIRCuz+JOm7Q0YT23MkZDUqvAwOYIx1FvedjJDRw6rk0Ry
oSr+/eKbb9P1/DzmRg6axAXVfSUYO2DRbUx6UztOkPkFwi/vD76q67ggyRpjRZ8UlwhAP5Jft/aS
hB04HJUvS5exQREJrdKEdCXpvYNldm0aXytGQqBNdqpDXROWHWtKKfv4Px7eA+xey8oVn8apIzEf
t2JcDDVFyq/wJtf6YEfhHSRXbgQgUYXdzqgGJz315Yrrpv0p6QDYdJW5P/IHvBdE/GAK5jkzeHDE
n1s6oaSYtCvxgZrGN/9H3/fbOS7UhawGII6jUwxLSwftrvfFgaHjtAqC7VmEvCaey8UI4o9wsVeA
EV5GVfW5AdapCTtxQbgAZTMAdlrQqTpBBp4xOLxX4G9nXVBZ9dkvs7VLxM9glPZcZ1HFqYskq0HI
cAfRINZ7Kb3xgN/3gCxqqlAIZpTrzySCbqb2Pxjjj1G8nbMYM3vQjr8mMoA4fEh181wUDYjsq6pg
NYWKjr3r1jMU6jx4r1pjp9Z40tJob44mImymhB7hCqqQre/r+Ahfzh1bR6PuNOrtd7BcaLntlUhT
FblEA0/tXdPwLmHAkmxeNbFSmxgQqiLpvcD/+lT/mCOOjXGibMGyG2SeKM3gjGHb0SQcbUW16UI0
vBOze0W5ln79+7b/wtYRnOeZgk6pQZ3jMDFwjO00AlUg9pHR0R5lSLUvv4oRiDjuvAYlhJGdC+rD
MAqbiUqnqCIX3YTe6hJ7Ol+aK/T5pax19UcCx1ReLt3UpPTYFau87yhRFGBXEHQth4Hf9YfiemnE
Iro6KIcaeP1qLqoglON5/HJ/YDe//K9OxloPRbQ1/RlgSItxUQBYeT0elV8aXd9sLVLWUXRYvehM
aXh+Bw9/SNFUwcTZZC/f9+r8BwNksVg+fLk6wbNKB+2Fzj48sO9MGl8za1VqTKaLS1Y7ZYHpcQgQ
CHmcINWprOBLETX1kpJwzN+hf9JGLBSWnsdiNxM0aKd2TUeIKFZGZaY7vbrVybmvtI0Qx6DcQ6gn
0u7QuHr8umetVgUPtEaGF+J19iTt3IGE155r1Wj1sUbhpVv5pbAZb8f8DGV5Ug6oyHrhcUVjgbsm
MOt89aLLfnzDN05WNp7STiA6jW6qAM64cCLZBubxbLiPmGbVQFEmD/c6HfsKxxdlm22iJ32tvIdr
H/7xohedWn+/+coJLsdRZDicS5HRKuRf05oIJ9XzguaD3CNtO4xRM6vOyRaBmE+pajaraOPwu3HP
3Nxt8ZTW3SaY8jUvv/uAHYFiqYla5wbDhxO/RUdzSRReNU6immpnXe3f1LzjqGXl87msREenkCPg
EokG9ridss2KWSkKO3ApphbRu2eGmDPs1cmzN5J1fjKXj4TjmeMiTeNCUQ6r6L9ySvfuCpI1X9ga
cmyylVeyVP5b6vGxjR2kpRkDGYAj50u2fUilJgRfWYQITr4pnSWtgW2SQSUZOzP4J+a9IX5e1amZ
7ix/AzlkhQTihuogWIt6UhGL41Ntms0dBO8dcrdFr1xOyGFsUA7Dd4nwn5OMEmjrBYhG9z0cH8lB
Uo+lgOmAkF8JMISP9v3PozoS/uzun66FJgR6ArLwoi1HCj8afqNjaBL0Whidk2wqbRUrxj6E/7XN
cASbza+LHk0MV6lfn4uiUx3w0KiH81f2D2QtKNbCpmXM2cCTcenZID1sZ/7YOdAeXlRwWzvRV4v3
j/8bosucNxa7tLrMiUMj7pCW5zThbYjuZonWMXfBcwNrhGQmqYtUT/5b46xj1uaTyKds+8bNS9xt
4MJhY8k5ciDHMhJ1VQ19X9y1sCZPc2M2+qPJA0V3nBj+PegGSRYUBt2UNW42SWkDgdImm2oalQxe
UNLiygCaCv3de/1vBzI54Py+6RzYs5LbYEok7ZUtxywXgaPKCja7sHKUuK8UAkjujJHpCL3sL2Pr
5S1Tidw5PijZnF2ndQDkMbgQb/rbp5HNKr17KP+eqG6iax6KYqG98VrWKLpDtbgATA+F3ctSscJc
s4SawmpJRCLMoyICfsBNnXyuRI1lIOjNf16bks9LfshB665hhXFQNPfIs2pbEVMMjQzX3rsIX6h8
/spEsvp5Y3AlcvDnpMrYBMYco4GUNQO5t0UcOG3id8lNdwTfHJUltqpE5EVNo6uY0IVr9DLV4XC0
vpoJvFnea0M3tWYCsabIsPyZ3Kl5JtCEM6xUaq936s51e+FtU74bdyuSU1/2/WRVhizw1HTOqURp
Ec/ThKelualc4Y9tptjHKGTfvtMvdslYlvPFMKI0Q/N0R6QcN6OTbT/JwbCSVwXGpY3PRj23X7Pa
Cc56ynoiIKIyqC0GjyhDFGFaEnkuGBKNbjrFtQ9+Ed5zxOkSivssk2R1ABN7xFvJGpJvJsWQDVB1
hHo9cO3TPn3j9fuHpIar7YlzNV8jhr/b78c5Je87JsKNmDhIYDOj6EQz86TxmGEbDHCZ3KzQwfOM
43XN34URn4tUW/4eU5gHTcRNqBMY9hZu+9tRcugRd2wKLwXeSNwu/E5G4YKymrFBeEcQs9ntmdGT
h9m5e4fIjeku46hJkcJ5fGv285sjbDXE5lOmmyfAcexU6OSJJaoYZvD7BKaw7zg/TQK98ouQj9yx
4zljYIxnuCTL/fp6A7uQ8usTEH/i0wSEIQqKo+QoMIMvIgXyiWrQ8cQB/QmFKCv3aGqjQ8ZhPNdY
QFka/Enli332RzIaz/gMaP+1SV4dVgsIZA5ekeQ399xRkS8pG91csuWYXArEzyb2fDvgcoCbYAtp
V5TKTEDIuZCm7Sv4L5pRPv6Dr9Jw+whu+gY3qVK+dpDzIn3FINql091pn/oCMYOKQARfbH+T9Owo
uxAvZghKiQ0fnAQ3E/5yrPLrHSPy3bqCwJUs26XZ5wconxa4U2KSKLlgDH0+4a2ELNCXMfPDdXvG
709IDN6yJz0zgZ1dTkGotKbGZFTXsI13DYFvbIk1uuRuR+uxv6TTeKPEPQYLw9FL3oWqNDt1bGZK
ZrqEwwPTLyuV37Y1h5Hy9Cl+32cHHCHWL+sSk2y+jSnULk2T699t4or38yOWoZuqMDv5AkTK7qCp
3GKPO4Sg6UhsMZ2O+7l6oayksYEm/J6wq+lb5FYcrCGBA5wA8Wn2IDwJlbaFu9B2+OjThtNBcybu
uoxR3ruT/sJaQbY7yXAD/h+pXzsER3le7FDGn/XKe2RuU6SBilyqy9+AdU181gYp+jRQrAmzkkAI
7e9D2qYB7f/VNNqBinql4HoC1XRM4Vo0z0y8BO7vn9/+56YwbVxW48r1CHDzFriQKsN5caiBPh3w
XMHGknrU+23TbnymPdbFBFY7E9+bwDtWhScwh/Xk/DFw8KS5yGdlYglHWGKf6QnkwSFP+e3Op2RF
gkJy2NsSnjiN1Frd33WDKjT73AfsSWGJwtmJZrGWoWmlOwL1f9tdzaJ2S1fxLu/GDJSW1Uo0SgMc
0AiNb2cCN8NxdWP0IcDoeQGZDBDYGHfLFJc/Zvbk49qn1bN4ZYx3OpgD69BmG6VZOP9Hp+GmCpWr
Wn5P2FZBiE0lH30QbJZZ/J5VSdu8Z9JH5tqEw/c8XXRTmTVHCcN+IE4y8qIM4VWsHEshPQgpZKB1
TtX3slgT0hyqnhR+UiB5TPoLzDGYWctrcs/2khFkLwK9/nOdEX5ln0ElzXk7TDoJNPpO8MkGDH+G
uGmfF63ilR7NkHwrjvKlyKFzc6bQJ8qgc9AM/GMT0u5Lzd6hkG1tVFeF3nM4Rg42no5VnnbIk/nW
2rG0lfM6rurW05BjfbGfitKWMK/fTxLO82mG7vDtKLPsbzIkt4xxikDYisdFe8pEo1PCno56ZYxq
7yZjMuicCLE/AKhsQX/8w0gheM8eLvVXjwQbmHe5rp8HqXH07i1oSqk7Emciw15I5HjCou6M0sKH
rKsP7LSaKRdjaYFS7QxMJmiFDNpBtw+6KjyFFLjOIArM9xgLER0lID4QVPWuBjw4p3uTGXppo5ln
8hNjNh3jEsvvbJaJQuOmDSSKzWV2sTVYqHZYd3QtXXrKhhWGms9MSBlhGbWobiSkPRoiqikWzg5k
BlyhBEn2fOt+/i0CKs51cSk1D3LRkaDIcccD7gxJ+u7xh9T2ve3pWqPUCOZcJSuAdoJHwm6EMCJN
5nRzU77zhcGlp74EwSYHsjFg0BydAJQEQVZul4stbDG79pUM94gU4Ujnwjni0fURxUDjawUCeiR1
vrI2qZ3kC2fTdJTlshc3RR+Z2ECLKDefo/bC22r/9VL8AH0CsOZdgS2rOATG88vjcdlY6qI5y1S+
pREcbA79WnaAt5iLu6/ggv5xorzYilqkhfCKlzxdJOR+PUbNjNbuwOvMTPq67pQPdZcZvYiaZ7Xm
+kI7wY6wrQ9UpsltbXDw6GzXCiyjQYtDKbrOTfszz2qvY5tR8j3FVpZou08P7xbdr6PlQT5Uh0oS
amSLiB8T5ARIW1IwCWxW6JIRNbFkHTvjAUghekGpFCNGnUELJbhsuB2fxJ0SNFD8Iyj8owtv675J
Ja+KMDwCUWNrPs7bpEOjKN0KVvr84sSIkkl+d9H0mg3hY9QlGz1JD4zV51wnvVQLJYnAZ8abDFPu
rYLlEHYM35wUg/TIVuPHfkWzmVq0rk0bA0Sw4wobTK8bm4UimL7RsHXd4GCTALYuWebE3Jpgjnhi
CBLx18y+2dRcm42y67zztl7lm5d3C9TIMzNds+Ff/hhE9ZuiP58e5A7NRxWOF5cYwkJ3b7QlYSoU
GvuwZ/UbRDy8YLV4l5FnoJGNvMdeSWK6nZ0wkRSQ+n0nGenJ2rTAK9xxj6rRg+xjyaoKx8UxpEgL
+8c0pNP/0Orfden21ov3fZB6AQusppnqWcKZcBE7Va0VSqIceKvTZTY4Y4glV2log7cqk2BVngs1
9MH9jyNGDh/cslHC79qTz6Jrwjtq7sTUsgPOOqKL2B6IXfmVGvIulVQzPhUrGPsPerDuBrMe0Ji+
1ZiXSXu5sAS3fYe5YiH/EqRJkUtPoCZLxi0lWGucStqgj1+yRfyp3+NJmXZhzsP1iz3jq9A/n58R
EGheWCpwU6yej2PWwjbg5kUYoHch/HPPzGC12EwPt9axWrgfVN6k4BNs1vk+vRkTl8OKnR2SC+hS
d5TsNa716lAZRQUY9xyhgm86/tVzKYGKOCxdd2rg90tV/z8TbAgAAq32RCrZmNpUFhZfG7G5CD5n
2Z7xGlJJjRqsgPkh2Th0kz7CBKhYlOd+KTVyph6wXMSqxBtMcTVV//o2EsY6tB+OgCR+6Kp6ZTyH
/Ppf90pWgLGHtOldWd5jiWFjvskU3ANBDQWAfTpDgxgGBv3Nbbf+ie4bi8CLJ7soVT9Nx/JlFp6m
ZapucKFziqljcOLm4M8D3CI/enPeldobnvd0VGos86qMXWEn/0rHN+ulIrCRcrb/lsZxLnvmTZ4f
FbGV9aS3WGkNOuNzu5lPhusv8eyn2Gw0i8WmjGHlvm6rvn7/P0F0ZGH8iDhHxuFCM7ATSfCvR+cm
b7fxEcDO5XDMlej4Ud3fleFh2tp2nmFAeH8czP8y7utMuJFJu+19ZgMIxRC21o//SCSwcALpNh5p
BvJZlOqvj9zpdpg8AKC2IuM324dQZTkdYVvIQ4Dxj6CmfxjZ4pQYDYLPYHXrLqpx+fAmY/GyO8gg
H/hZ2SsPHGGqHqDqFHluOC3U67Bo1PfBKUIc6lCMWhr3N8Osq0s+JuwRo1IIm4/gQc4uOEgMhOKc
jiaJupsve7K96Ye07R6zzZo/d38jdonc/K77vTbx5Y25w2wCjD3AK7A6KHvbwQm+FoWYI+DsYrCh
6wPxLA1xDN4MaOUuzyZrTRaiKQbnQwQKodcbsEWyuH/gNRFQl+9TuPhiGeSXodLoQFsKyeY0sqZ2
KF1Lbucbi20FvPKo8Pl/YRY02hXCLhYdbSCUOo+3mGqRH/GCabXIsYXAT7aTdhcVEPUCm8LK91Ov
yteJoJ+Ekrwcq32XdZWDn216reHPKcPO0Wf+aVvkLoEeePP6NXh/HPBLwLp2sVbY/h/i9rMUk4XS
DoEc3oxK31VyNF+0oNptkzqr7UKoTAeUyHJd0fywPOrAmPDyuhiidk3upXYdXd9dh/2/g2F7uncS
NgZyUrPF2ywT1h7eXJtqz3sNHgF2jaZym7FZmqSK7fInbkaIA6o7VV/bdQCJnyGIEWpjyogPokRF
HR9MoIu8zSDVNOvDToWkJ8r8Btk7Th1kr6nLnhKsaWH51R0RPV6KknVOXoEQLia93DSwDBlazaEd
2BPdLv5b9hYenbyzIYb6mx9PnN45z3CS18EExqNiElmDcb0qs8gN8l9YNWLVlK84tixB2JjpkQEZ
jNTtWhwdlKnQ0Cwu8Svgs1QfTQ98Rx31hAG1jDmUrp+ElFP60NoxsEKfJAdoI8jSL9PJPevNbHkI
znFtItEU55Nf11ZGg9FVN50HyspLpkEc9iE1kq4P6elEF9d0ma8SyVLV8OLPKU9TpZYuYwqjrWiW
kVobI5WjaIFTScMSNR5TPPgvyUYxtOPdZkwChjwGN5gOQ55qYEu81wmtA1iV7jeQbCHB0+AGQYZH
GLJWHl4+oRzFhyH3NFfUgl/H6IhEvvHG8Gd6psUmPrSKIyz/jbGTip+ihr6lG6W282ZhfmSuBwhr
s6MVgsLju8/mCMUlTeCcjZHJ5AxGh9qc0bnjGwSiiaucVdC2LaDufOCix98Qj2dwieEzIMLe40gr
RWU4EyM/JgWu1t/YyXmyxbww3HBgA9jBVvYeW/6RvfhRyJRvjxJten67PqSW4aeOwEFzDPDr3631
69GOgk5sWIAQM7VtcKHABz4dcSXe3yCcWYeCXMqvXK804pX+uaEr3rxxPhpnjDH7j0xx/4ayy6gV
IAAVoA+hR+1AbNi2mUIUgxpmECqMp37YFdMTfN2Q2zCOZlNKIxazHW2dmIphFlQjlY6MbCdL/YNY
BeZJDlXuCLz8QaLRtzl5NkdVLC4ERLQClO+6l6VX54xB8kk5YEEtByzH9MD9vEMDGeq6Hg39IPAC
CKcXf1/KvZlpxRfzjL6IcU9UW+DP8V9jsx89zB0WyZJnXMO4v+6snRrMJj5P5m848cHMxXqkcbVK
pPQtnIXJiQxbLPA+bUdJMBHpZBLEHtCGsBqGfcOABPv/X0BkWQ7JKLFrPXlW2HMDM3GMD4LAeFGj
9yA3XcOtocgFbZ4Bjw27+5r0Nby1F7MQXf6KNbRmfIsTcX+NFYoA1hSNpSBhfFGhsj1Wqs2Fx8G5
c/AWTVJ2TqUin1fX+8lsITI68R1JmSQrYUPQFXTx+ZMWy+wNmK/9RGvbx+Hud1oIUIwbwyr3vvMc
VfG06GLxG3iO7qLjOyvDEtIsdTHxs5LMbvA8/hwYKTXDKKx0WHgT1FqoLx3Wa583HpSXIrFDluwQ
hYsD+5nu6RV1m0dBHuHPGTXbe5MWgVVx1osOEaogTV4OO9ITv/Fnp+yA7mTw/77NJkyEq/R2Pzuz
SrCeUFNtVY05sMHFhJm+shayhZZCxLtePLQoSKdnY42wBlfjQo2OZXEh0BE18Cm/2intyuHmrQ8w
aWgav+rJ4/xY12OiHN/WIRq4nwNnq2mXd1/+AwyqWko9+KUZY3GHzJ6VO7kPDZdbfKW3EDvnmvDa
CcVwd2WWpKeMyQJoV1XbcpjMqApQuF5IOkzgscBKmyGYUvE8vYC/APaHJF1nd/m4Yl1LtRo8sVSE
YnWv2DRmNbY3KV/ggsdyESA6BGcN3wDFPXJPtyR5Hok9eHdhDIhnfDS9XydPHkPuw+dd1kiICuLh
V5Wt6owIVPL3GaY4zXn+OWx/mB0ZELISzxATLb1HZyGGMudjqB4Sy1vmagB41dSB7izBdGfzLhAZ
m7PiURolAr5qIZOvwEovoOwvX8bg4x/KU8AYJ6pBGQde6ehWry0mSRRVN1QtxJnw3u9EDDk0D8DU
gWjknnb2Ivg16nvjTPJ9TzyxsjyLYv0F+kAHHZwwA94c7NVcMJMSP22GNemlkLGYxwcS1AZYSt6H
j5Wa01G/n4MfaiZNI6WcO/Mj905Ljg3wO7Ew7EM3YGEuH1AIKHk2ywNSQPJ8YgoH1iWBQCQI1+xj
YphjUyuXybsZ5okX/GCsrxP1cCg08MdK0pkPvY/CFHxUC+XnrkjXLZqNDEP60Ef3631gpUeAXfNw
bbnbSDdaYHN/UvwsJjaFjbhdpSc1ClfdEsFcp/WjQjwyNxKds5MkbaSMHcZuyj8jENbgLzIn9tAe
pm7yWvnx7RoiRiD4PckquNLmIroWwxNjo9B4osBn+nZnOa90lWGzLqMKlTRmFLSh4K8DKeCDEFYh
M/Zyfb7GDZUOs7KhPB3SI45dec84oU5eMSYtVYwzZxhKVC19EfgiTU0ySNdH+amIEYyszBMruTRa
Nq9kMhKxEVZSpOuYFzxK2+mwkLfQiAYs/AwsGQVfnA1GfLW5o7rMD+WXkQVolmx8dxadQ5z3SF65
FoaDVpB6CJ//sfd8I4JaVk+XyX6gOWjphT69hWQqHnN7sjv8m1xYC+XbjNSmw3FwjiBsi4Outnqd
cvllL2PMbq9sOHtO6wUUMl8MV8kQgLJFvWN197yrI/I7AZ8QWsR83KP+quHG5fyr5fguiDTp1zl1
AbSYQfaV/r0VL/mqQBJuOfbqlvvBT76htGcqeCndrCoI1O/9O1mEUp9XikXg5gz4eT47GQ1eZe0Q
KVZ5lyPKffk/xZGco3QTe9gQIuHwx0sbWsOP2vS7i8UvlsvaYm6f/AJ+fXsRXA1HfdgPm7Jy9Lhj
T2V9yTkWinY/SvLCCogGbLK+OCOgClL/gJU76u9IxTNCM98UrGYOaCc+3KEW6gOfbe3WOhbLXU4O
pgbiN1mFFQhKd76wPnpS2CzsTBA4SYAVXgg/ycHxipgEPOPs/uXYmeBs2Aq117TlkBqU0PUyO172
vrlHld7V+b+qOLeqTzuzUHr8NkcPqR/khVz3DW/v56vKoHTQpBf3LxIAfB1skNTDUQJA3+IAFgi8
1GVubu5VEtRK7hwbzUdOPwfG5oGqJkLik3Ci+dDEFA/CQW83CZW6jmbJ/gifssZ07o4hebmwFqet
SP7YFq13XGBmFY8cxnkANEaYVfqSFiXiYwwCaWbLaezPpq96qVillps8349OXLm+nb3aRN098n9d
uaPr8cUdWvwv8YvfCAKX1vtA6qnVk53ptN7Jlf1PeGGd0CQig6nnXn4g+SrUMgwqYpsHTBuj1KfN
Su9BsutoR959VGvP5f8SgnQB7k2UXw79WdLsm1QA1awGvVDlL5raPdDkX05mwnJVy+zLubk7PJlH
vXe4m8J9MVqtudCE7aafvIik2SBrIuitWzChQ9O6O5PiI6zGir9h7QV/Uq4QD+Y25toBedY8Dmgz
Oj5gFB2pZqZKVtnIACxXOXUhvaUyUELsNHwIHYNMap3j34dGFy06/3LyWAW26cRtVJwE95lflwxu
MVs5dmNMZcVscj2iUGiFXQELnl8HW2hNZJfBQozJ5th0S/c/xdy4xabdB1g3zm/5hF8REIBWRxs1
VWi4HIgeY1ffItFGJ/E6W5eIlo663Dtgc0evijCbH0FGx7i1EPWwnFN6bOV8UuxNYRVp4TJN/iSD
HAki9DqJO/8kBaTS5Kfffz60q1BFY1MlOQX9PsSosT4HFPkVYZm8hkA0iaeG/wehnNbLJc7N3xc3
4Em3Mv8ZPn96cvkiUrunV9hH2TDv5smyuQp4IrwfHhdMyjCvNQI55uJiYgvvTrEbw91msbgblWmb
hnQtx0Ug7XSC3qbOqTU75B7zCv1d+PdFjPipFSS4sGxB6LyAa4cLbNOOs6K9nj/3jL5BkczS/35o
YIJ/1G8jbEmkmC2j04n/UiU/WWrfoMbSGNmFflxN1oonI2ul+LCm5dnUCNmcxmC0BFKbYUuwQh5P
4EXKShS7LX/aQARHl/GZqofeNnvcLoEmzmK1ngdb0W+Eo1HWIqwXFZ+7SOXNws4B9vsNXmZzGKFp
2FxF897G0Xu+1Zn0IMUnxutKKQ0tauc0i8EUqAauJ57AwITM7e+pzz1jbhz3PeYMj1wvG8RPEeY2
HT7EgYGh7Wp+ImnOZrG8YLcldYACPsPibs+MJOfyhZEfM8YjUfG+h2yKjKaX0sa1HIPaK3iLzznh
sgdcUqezyVK0tzcoZIABFwYA0F6oTx7ykx+FDUiHIXCst1lZlOEEtAPjFqFaaBbO7D0OD96MMfqI
pxiRJMJLaXGoZFIo+aMkBF7VI60VuU2N9ru7dO6PU44d3sbn4X/o1n2yKxQko2svp5BhLKIBJbvh
GMBX63RIGPB59itSXm30FzGeWS5y4We4DZ9689JYTOmt4AeCZIC1zOoZN6iXZHprk64J4t4ULIEu
BkdWoKE7PZg+6HnOumazTV9eUBpQjPIsF4B1hJfnOc/joFZfrnAo1b1zsL53k2/fcRog9T/MzOM+
ukOpDL1mALppMDeeaDy0/wRd4YOA+exRY7VC6P2FClgMl3Z4KU+E669BnxakP00TktPDhGHobuH/
vfayAoGYCwvd9GV/FpqZVk0E4tVAG9e26VeWPcDbL18zWMGfUilkk4HbK2jSsljuSpSfcWyuzfDY
fbwGVt20wH+T8EBVWqcDMwxoRPUucTaKTGNWzfc1fSEEGdgJgMvaJWU051zMtdjGcq2bCNNWxsBY
Js07PCM6iN3AivACpDa68zQLuxG6fMys7ioU2r2cb5POrKN0OE4M8uF9Dqt8bo4qQBrQBHoCGkEc
WflJegPunDB0WEsA4wZzV+e7lHfga5UcXTyTIqnuxphcdoBFVb0HeAKdhrgdJ3twUhvhMzw/HT6N
fIyQTiL9ipj7bAx0xxurB5RdmPDvYVe0iOkSsGGcPVvbe3dXLcSR+xcqP74Vn9OR9kFCv7KkTFcv
hDEMD5aI0hzKnuNdOyR0hokmwSO61UEggN4GH+P128wW8Cuoln8hjpkRV2CC8r0/sv/f86aUgkGh
BgDT/y86HIyjscs6nSvc/993pJBBrQCb2B/w7mXYBmC2ETK+dfvscZcWvVzAUhFoKa7hSnrNH5Sm
zn9ANOE2jlInAHbweASyCMh+nEpkp4Ir5X+cDM14TL+1c47v5XIizRyQc1J++6sbp3Yr75lF313j
tJAHTSY62r/7g1W8q2MSHrwcMiMwwGdilpJr7m4CZq4R3kvYeKJFOFlGrkl3uYtodIDUD7KNs37o
2SHdktn8+WGleuXvrqII47J/IbSjx3II1ZUH0pweHZmkLW9Ifr4FpaC0wJBiIlltbRjGDNgjY6d0
OP7FD5mGYmq5xc9QgQLSL5RF9+CNwq4XjCOtdmAYezYypLx7foAgWJRrSY5lrrc9Qhkc7iZ6bfu3
Kr3iVzZBKa/baQHTdsF3NqnxP/7BhpAJ8BO6YCufmytlfb0Kal/cHCJJQhaQOumcGia4g28vxhVD
wMmIgWdLQRV3qxTENa3tT2QMw0Hl91hsPGQfk6zDEZuR0AsttkoB5AhLkpDf1ps5P7jS9IJ+su1O
GgVl7TIL2gmmRy9Hyp0Khnx6/qWEAwarzfZdJJlXCXg1sXIQNcAE9mnW14/0Se0OaejgTLLQk5yw
j10sAvpOQxwyrYjir21DFwd9epT8IyCAPARxssPdhg6EuLocvHLGJ8AXl5xVC6GjDMw1M0/2Ba9F
NIL773CEDYyCXB9AVM1JPekYHiwixFzIi5bEOoi7I0QcQ+q+kQ1pKUvDuG5YpsiTrEuL4X8/nYLU
wr9qJi2u9/fFcyA+T7+iKm6k0q6G9bW/3cscg53fHaYC6SWcJMeF1QXOIml5Fy4mYN0oCMolBAcn
iMRLLbMFwReBY7tTEjHHWu/CB19fgCtmrJ/eWSpjXYKIdprDUZ9FRnQJT4TYN9hWBDr/V1/02YBb
TkL5S5cX1lqgAFMAHwmv1pnKA+UO5iZcXsLWxC21idkeDYku9Pmn93fx1rCb2Uj6FfLj+5lCseO/
L91CleVGh5cJiwILziET2Uk3aN+ukrcOj7VHMNmkULK+l2SZI5YbhRIDdVOLGcPsZkRlpXBlUjFL
/UXPC2Zw+KVLZ4YoyrPUkDLrgPioLBNXkaNGo35DASRr1JqMZwBzNKA2HCOqyc27soDNyeBHQghS
zuKCshU56oxyRQNveHZdmGWuVMr8xbcOqqSaJWXyh7jektWeI10ttiwDiCnXhNtSKnc/z/bDC39o
9bUWKUVDwOmJuoxoMEqRxjoTmZY1Y5g5h/uDJqUtcbFYfd8HXbCzOTZDvaa29SWiD+YkKILjpBPG
xwd1RnFaUTeCOSAhmUPnSr5gjP8CfAN14nNO+oHmmFa19+f2QFV1+eq1ghWd3odlg51MyDMASITu
51Xc+e6le50uK5Nj4tNIcqnS+a1sBC8p9XCQPe6aU13UNTDo8eXNfFhjjMUKjlpTXKUk8S0Ipql2
HlwHLIVHb4WCoj9wX4+Qzl7nF3CsChN4uA5ATQ9Mn6oKIGl/o8LErAEBMBX6ptdns/Q9n0TNVTnm
BpzVKmxwK4K7JUZDBWOmCR81lWgD+ynOmnjyyAd8osAQDpQmj7u8us+gR2hKK1llta1d3IZ5uFI7
8bNuzkcimLriSJ9PQqQAJYRsnfdw+g7/3QAwm117qHpRDpX8YN6eybNSWtQnHBM4rNsj1wo1wSyK
z4+UhG0h3OIpc+xM21naZUYG/p6uOmd5OK7VewcNu4Edf9b3VlgjQktsRfKpnwAgNdfVz/PbG+29
ws89aFZTxUAV2qV1N/xUrgWVoJoJN6nnenDoXNxXyVZwBwWXdnW94i2mUUYhYrif8C8bSBn/b1Fa
CgQeOB4URI2xU4iZVU9izT3ZYXagDv0MOcop0gMh3D5payjnS4DpcU8CCYhjU9Id4AWZoaP492d6
SJF1nOnSINs0FarQrXPowM/PWjprGzpoUgy31uHtkeogHICU82ZT6iMI1iBv8ROdvWXg1C79stIQ
XS1J0fIJHo37gbA1ClTSe1SzaP537Jf/NOnNCmDYuHJ3aOGUMXJsT0JArrWS7TWpA47TXj5urL5P
2V7M4rz4JzLOp5dQyfcr8Ird2hLk6LpVvxPyLK4M7PBxmRyKE23aPXQZ2R5mdOKyAn/PKJxSNROE
YRUsVMWKVtjVyWSiwT8t4QE6Jh3HuveKpiX5oWsHlOjsqqbnBH/VleME4Vgxx0laRt/gN8zoy7cy
nQ8PRD4lpD5lcNtIYTtufpF4iQ3Z82s58ty/nBWIBIthST0+6TxcIK0m6/sw/NaoY5odixnpYeWS
pEpV/+wYyjUDYuaC1PveAQSujtJWuYhlbaicsChOdPLTImFmh51TcrrvtooGlkidizt8vp4SHGci
Ry3bqxLqzlwVPrcg9b4S5yPVDUD1yDTE8A6AFVLLGwoGyxCZKK0vShVuWX8kOdpUOspjduoF+g/5
3QCfD+2BdkcfTKr/OQm1j37QVhfTarWF5/ubNRbf/t8jz85U7JNdD1zSoKEMqA5XwRTJ0hKutZ+T
slEiVmJZ+Zli4wVxQjK8KiqcabASBlZsQPygkeuM/H5/deEtq+rV0G2P9ORnxeNTEsbzolxbZXD1
OLuNVXIiyVWt/pC9/uoY/nYJdPbOPBbNh1Ky6a27JtikREnkIaUUCr6BMnQWDHkP/DY4/ECISJFB
Fs8pDzGFDKHpP01KOgv6lclBOOMcsTWY1pSEtEAv9Ao/lEBxdAbg5NmX31WhGSyXTV/bYi2almeN
2obduybqUkNER2GpmMSCocX2KqUJRV2J0UAKQiwmmSJdAyNRNvs2cf0EwHLu5r5wwcQDU5TIYvW7
rBxjvDsPYVtSEJvR+8qctLLj2U8mwCw18l7y2/BfKQ0fqz9G59rZMk9mj2YDZtdfmrbIzzSgfL83
wc3ZcH69RvFUwDFn3jjgK6Nzb5cHO3vQfCRd5vs7q2XJsgrlvKCaSY39tXhT9wNa+eTlIc2hNRn9
IqQz834KumosiZs2wmIeHPwNBT9CLK2rJDUrm6/3w4y8WvCrYLZnoRYTx4W0JjDKM1KPYkCoeYIu
PfpRkRq/OeeRaegzCPBAzwRYsmPKYni1s/OyjQudpU8sH1acEJ7qEQwgqI/6347JWACNBWguvFgx
R/jCHj/Y2pLNm1em3bVOKhtazQEIxbp2zG/zxLCHCk/Bh6c7c59wI7N8TaQ9OgtzSIzEGmEG9oQ8
1+o8azjsF4wrxMwSn/K90+wGR4uNkv9/O/kr5iBoWO7ajh3TGvjZIeP07/newojy8sFDyIDk3Zs0
LZ0gPOOgLBtKHR0aMILC2oUFEelV9uvHt8cY0828xbhtYoxy1ZXhF7F0X8htp6e4nUpV7lWrALE8
xlitKFTAAhuj1cfhK5/56sqUcNZYgaQNTNG3NxiBpKuUoWnECfYyiJGhLzALl0bmbuditIQ3borv
pvcudh2PG6LE7Le4TgHDh/1gz1Jo7z9dHcfIyJ3JF66i13cvH5/3zelFTAI5+scOj978FOyhRZ4x
w376D+Cpwl79O9ewlFbb/g0B+1Xi6DUY+eJWkMhLsDyeW1gzr/fIANNlEYxAqCu9ytf5rbeL9U5+
KoQOG2A/GTWBX/vrcsPSZK/XaPzX26aHSt/le1XR46bLVjR36NMpcOrSlwVUDCQ/F8wX2Nd1l2Oq
+h8HEaJGuuUo+0L828H+BPWUxz8Nsa7D8JY0NVmE5Cjvh0XBoeI236z9EuZNVQtRPFb3xPU7IP55
Ahk8DaSu/SHBgiegLDPFnLQjgw4fsJA8FiU9Z69LkGUwTj1EGYN94sbUcGxI9Z8Z1YFLGqMoSZLC
SnGc4Ak0yMUl6apWgfP9Wa2QydN06Z3GrfCRn7nASYtLjp47hVhksX9CGFP/Ic+v7h3acQpAQHpA
2SWnwNQfBX3jPRquOCmrd2Cq08mgOQCGAoG8zhIH40A85G0ZM3ta7DfZ5Tzz8VOdl2mZD/hJXOKj
JLr6nyPA8t0LvRKNuxqjw1yYkeeC6ApVc6BHzLy8FIJd52WzECetMcz+pgW5otWcG20UrDsgKRI6
ZkEd5/wdJIZKVxgcSWMSMTZ5iAtvQmSpJdRf5f9u0E2dZbUxzWweT95y4oL8atQBEHs1izDGWhi9
EaK2F+Wm2HxwST5LPvAUzIYIOhjZ0a5fUo58H3odgqY9QB+jnMPRNKeAMSDlZNd0iai3B9CZperx
2PfvkWfxpjK2FnDO+b0gba6DvRVk8YdTUJL+MO7Oeds7vsRDbTlYiB0WWCqqUqc9Du1NQIotCr1I
PUArSDp3cYf121btfFMeE/x3x3eIROk5Sj0IgBHKvwCpuX4Zepd/wXqztvJUO8d8IZncRhHwZ9H/
PLQ6Nd9mxGJoMoEQrtAmy2Na5QB+Z5lUnRwtfr/cBM+Gc0XgbMmEwoiJB2z9aHenNcvSHHPDywwK
KA+bejApYre+UVbQYcFnxgDVKYWm6yP4ULYKfTFiHkYxZJWEAfKHjwUjmD9/zBamRGiQ07qRs4dH
5hcoWhlRhPkt2CA+KLKTIdBtS1PD0VO1HnMogy6iubYErAI11D6Eyt8TMZN7xWb1r3B1fqJ3umpD
+u6+wXhNuxveX6bzWs9RT9IGp8OfVHr9cnUV4M1uPaEjanpeVibU3tcZXbBk3V4j1iptnAK+Knrq
0lO2W4W5/WByBOmrGoEU2PlycHaoL0denxKHXaPJQRTxK5+me386mkGMjoRX7SUXxISkUdIolfZb
SHrP/zRJXVbYXkf18Vudc38IqUMp8l6uBYzKYmCm6pthBIAqtm5373Y4tsO+iw9RaVU87YKCMMgc
D63tg10UfPV3463QvUjicEqQuFvhfUxrEwzB4tI/9E/LoaeK3eiXR4tS4+uvxDq5gMa7q2ZT/TxB
KN8srgYtgxiQzZBHofTWTC2LKWNyan89mnHVTisq/1oq8jzASu+y3pXOrFdsUlr+DmrXLwbQy4Hm
4ptthl8jwrXjXqEnqOCAFrBEeAGQoAkErEAKxHTE4UrXODK/A63Hz/afNhNKLCEdYoZ9TPt91yl/
1VL1t+VE0bcdMJEl4oe9BsRTqUYjLMult/I7U+qjjgxs4+JEmJEFYjHVKPv5wL95u6zhqvEXq2mk
D5QoNCbnGcFWFlRmTv0Kuvv3jST5y+S/6wDp6RLW/mA/0t3bf1gRnvrHfzYS1npLVfdI7Jv60YHS
y/vYiplbYDnN8P6FCDOdYgS5Cs9AYTadYH07q06zCbsALj3SCuh/PeC2BN0vuTOpdkrN2OEBTpfD
FbhQ+7MPxgbXkSMpMDRxx5MbXjAmUWWsI025Lp3vkwT+5jQP8WmW3kSm5Ut5bJ9PtUDSwJSDCTrI
Qx60ai3W4TFWrnOixVocRXC0d1BU1fhq4tz6I5huHFmjSg/xpl50AcR9YZYodXCYeKlILfkLglGM
et79MUKqEtNCKd4FSnk9v2iqNCxSZcSGOhQJWiPI8hecvYU1kUCsOFJfK+2kh/8yPqhY+J2eyZ75
Mln9Qa+dgOmkfhtSMyVmeTlKA4WHO/jhN2svQw0m9EUUsjvwZ/fFiMkD7AzH1ex4hjrFYf717+H7
eWFFrnOuQhx9HahLsJw8gRj3XKF8XqXjqzLs1iTABOiubIgKjLHLRJuteGmNGk1LUBmsoYnBjg7B
ONJMOs9enRGi97mnuuGJe81KUZVp6qwAATbQKmmtB84KXkJFcnzXqx0TWrmSieLYkyB3sHHmrUPL
W3uqFFIrL6skjAp8cMtB9s0xZkhx+cjHRp9PpJ+C/0vuYf+KrAtP8KwB7BvbXQaStbr00W4KGMCr
LIJwqNU/whT+kxFLWEFomALPEkWbeazdUlIUdgBm/YN13kYjNAA57dhNznpLPnRnQPexWE7JAtMr
3SbQWRBxJf+b7NPwBFvW4uf16LR7DcNNk1GOfoDwIyFDoP4B03tZZzH1Ku1kInmVPn6qJPpFMz2A
5Dz8y50txQ173IN003KD4+c+x2+Rakex5nnbXJNEZXJUfHcKQGM0Sj/6ilFGbrZp6Q9s1JUJ88a2
8ecsGxAFepFTpOtUQnpOW3U6/UDen/IP9mCPJJ1JnEGLfA9zzez2ucca9vppMEmD+p66ZcFOcdcN
s5vak2pZzx1zIYuJMZQ/amjhSzStF5NX/ztnBJAcVjGFg1mf+QO3SWyGDC6DkHsRnoy08jj0IMEK
8SH+LMpcpS6ofFFbinX9R1O2SV4Jfk9d4B5QaGrf8xJ7LilnhpU1QUZqNeEJ6JYIDUwTzEvS383y
ZF2aLMKXJaTYLpe4U6Sh41w2+VeyRUhmp8GfCdpK6pDv6c0aSMOoWnPtYbv57cXCDxQB+h5JRZtn
8O0LIYjEz9vHQkX5mDX3t1FVR1myhCeMB7xDRLQ59h+eSI4/rjKGkTvbeYQMGposdBkdoP3PJ4zb
hzO6r1V9fnbu5Ev+ZpyV+nMBnY5zedPtyNDDq5QAYYha2TRL87C9f77tWJQaQK6U4lcgyNILljH6
tgw1f95n6trTi5tLjqbq8NPMv988sOyxIQ43rJ1zUuH0khU7gzY4EqpqXDI2niDt/8f084cCZIxZ
m1cBICGuGObHFh/aE4pxddWNYpxUE13a8toIQkKWQ62pjYVM18Y8kudT9oZ9W7MTcpTs5ifLRP+l
CYZgF5kzpWxafGef4gtEswmLVWksN+Gv9I7OdaaCrdu2HvCAkv0A5aS/otIo5MyEp30PXf7touRg
eBtzbZaRhsBBBtVkLtDGgrffUFAD0ZDL9X43mhuCgnls5QiQ4xZumjBPSxQpo8m+s7njpK8qPcDB
tLevpWhgCWqDgjl0vblP2DFSZUQS/CLjdAY/7ZQQkeVjCN17ZQN4drTBBjJmr4RzpN+Oe6tv8epG
FAUpXPHXYttZDj5B1bk/fNQP5uaoy3bV+16xYGy1Mp/l8+y0dxiWVZDTQC/MrGPDWpm5Sw4du8VR
V9iirLICDE4XAWP2yf+54KkUkWUbefHNsK2XnoYOXEu/IKQE92yD3oQPFaECiZ2SxdcLqaAljsAa
kwVjpBt/r78RtBncv3E9iC0mkkGH66q9zoqwmmN/c6bZPFZlgYfXaU/X3L9svFw3AqnD1tJr8rDe
ro2A2nP6VrGy2TfezE+zp09KKrccyqcY6UbHCn3IJXzJFHUyq6A8susiWNJFr/gb5CztUtUrYK3E
b0Z5acPIlCmhFw3e2rbXpHeBNG40GJb1NXuDJZSsK+2Zjpww/YiolPMTvAY8jSXKD3+HL4Jgj9X+
LIwpjRo9OsLu9chpbiK9lXYLEAw9PPo/CA8t361DxpAbPheVA/sZpVCgMVdBJuHv/5RZ0O6KP/Tc
atLeDllET0Dd0SPwZmhw4pUvJ3enk3TO5bpjIyNk8Kena9ayDUuJTMSMGC6RBrrNGrLVJ3/nc9Vx
cjdP/Euc6PhJSrPOyWk9peRd4Di7UgwqGeFb+NjQJEugUxS0ug+qdnocDWGMsxFupan34WOK0X+U
tq9n13PPMgxDfva7SD/3iDMApute1/nlogVdKEmyUdfU31wMAdkiSokYI4YheagrfZ7nihoIa3C/
k96uGa9nbO5VsZqbLynyrmGQiLt03P5aca5i8NwIBAdzgTMOi8wkXuWkjZuEn1DLXPc5T8jGMWw7
BpDj5l+w38ZblCjqewDjuUR+DujWGFM3IvOBMm+aqaQXIBORJp+IycRIcuxZLY+M2SRNe/yWJCJJ
qsPa3OWyNDl2lAi2oH5EVGHU+PEAr8MYtMHdAUrq8qkHqlUSHRSuEnjMSCzthzu7osQYyx+ll6hX
vOBpiiiE8R3ddfI8trOkyQs9QIid5RoWP2fg7UDGOce9sr9W1HSPfl6hIu6ImGAWvqOHbfs/3jCk
iyESqTCNai7rS96cNI2mQzNy0oOmKsaU65SMrYkWwqaqFIXBbxucmWd40d90rYRcoCZzEhmurOX0
2G/Psn+DI9PWgr8P8I5ya4djS0Vf7VSuUgFQZdB2o/No9HaGyoUrx7z92fkfgFx8LTZH6k9C1Y70
ejaKzuEKFsLa6nHcvoX9T7v+HXlyR1OgVhoJkgXVuyec0gGk4DMWCU2/Qos2jyqNyjXMS14mQ/sc
4ay/doHhLo2g1Q5x7Wqn2t+k+non1DUrtRf4wgseAKbH2A8Eak7/9Ci5mIa1BeIS2k9zBvKiuKp2
aXPSPT/an5JqB9OvhITvu0cCESBvVpROfMGkE3igVt2oZ7gmAj+2VGM/bXbBC/AwA8qoVZVv+vY1
EF+jSR4L/kosbUGmSu2poig2tbIq+BSIzPuMAdf9treurn/vzHiyKXQkPqvOIoUNcQ72BazodX/q
KD+KoG5c6nruuYQlzAiaJH798g1KiPbq1OxS5xMX6cuGlgCGvNoj4wk/fOiHwUEhg7dwBEqhEjZL
DmTxzKn5JmqOoDfECuStjJFuOXnvRl4E+/nna0Rf83aTivAmjnXOqTdIhJR/ucIB1zkcjXJbQZVL
HW0bn4SUJlMGov4kuD1S+33+MHRmmFh4InAYvVIoF6Y7NF9G5se6tUsGGS5RF4hBsOzmCstcn11D
rMPUgEuny113lOHqFh8sUgW3DjuDsO7ZSEZBa2TlbwSF+ztse7QDFjOtSFhqLUTG5uFmJOzOQefr
CxMBAPnHs9Q11cDCr1lbmb+w72dSjYuzR6EpBPuUQ+bPYLjQHS99YayqHVA+5HhLJQ48UtTK3kwd
W6LFB7256z6h4odT71xzZmwVyuuo7gX/baIycF28wTj7UGq/FBttoEGIOEd4WBZF9qKNYWaQNlyY
jAYhvi/PrzOtbwUirDuaClTE0w5F2DvFZ+Ue/AGeBnMN2cNfBZBeyLjWmu4YgY5DzX5jfxr3uONE
WwONQBRx/MldhyyaU9OYkwox54VeB6AfjU5H7ebUgyJoQptVZ8+oDEZ/Uc5VLbKgi3KSjYgtv0Vx
5akMbce74o32z5XjvtulOtAKhg8PtzHqmeDX/Z0uUozMvLnC0BfCRuUNRfAum33/IL1nHsb5GT8R
DdQ8yGN33Cm0+f7DWPXXamYHzwmnRAf3+hu/J/1AdkC2d8Fl3LF8czQDm13rkzYYugtak8uiYvp8
LExp6SYZfgj+AUbLaHS/7skRFIwYn4CFcIFi7kISeYaqvSFTbBv+PCDPNpafIytEtO54dYenEenL
vGbrqRU7TSPb6LOBTE0KrRmp9c1iKI5s925t4wZ59wFAy/ZyTyBH6ep4XdInG14wB7nyuXectZ4Q
pKfH6FgSJUBRCbzliogBEiPXVslD9p2SXypYfJuZMoCm5zWpAszB24VEvATK6pLP4qhp854Bas8C
XLeXbAC8NwCH+ZSHKGQpEUWRW1URnU80yjt42xyYMEugTm7B78mec/bJ3zRsjFQ2Ewv2qPYD/JDo
0ETgsN3dP6N5MpzxG3huYQaFQh4SU19DwdrTSDLLCITTywpsdEBxwBIl2izv2+fvXAlLCsZSDRpr
mKJyqqnKerVjhmnRR/ABF7/8uzlVrxly5ghreleQT/w4MmFFrowHVU2N4Pj2F0tuCmyH+mjmzpLs
Eq7Ta4UL7BNXVRsR0m3BZSznW+LKnH+63t7yEXXsofZjTXoQbMg4qNqGNkgel90PURAEuAQmSa8q
2CAlCXJim5EPoaTEepxHTHxhvjxoiorRhoDt5qnCSQ4UzH6n0ehVoziH76u4Q4q58jg4rHFKbfGX
Vd10CJTo3qUf/aD+b++nuZ4EvCzdSj9wi9BO9Gq63NEctu0/s0TMpbxh9G4xwjDGWbKm5Zb2z6Lh
+b8b9W2GpCSj0cimlg187BqoXwXFD6DmW86/QF+sU/eVe/L2oZMK/qFz4fow0a+F/LVe5QgXpp17
Hc99jcc963FrgOdE4A2WH7KZVebIeyotw78DKtg/xE4SzBJiHzRSUDzmlJo3Lqb7e66DxaLyZO3N
e1DUY4qzYWIotazdMbmJKZbE3kqMSimMJfSDwOT86iuGNd1IdZkkUlnKE5Jxd/WSsGl2HuKfMlqG
5nyUvOS15lbWArm31kN1GY7uLPJNQkYVXJLYff5mv7mTknLUSHNNaiR8QK8HAxq6PP0IvrVv48Q6
3ZnF/1FZIItxWC0ol2MxoAq6DIR11N90wsaSLPUzPgvf392R8+Ji6F/xCgSA9z+2653Fl2qhZbYT
vcNX+107pbwhxmKpB1oCtNiN4l/ID6KHIjNp+Y7m8YxN4J+U5L9nH6KR+9ux1/JQwNffnYD46ftg
ZMcBuKA5SuiwizYBn0+a80GXAEbZn269pRfl+vIyogmpJqaJbFmc9kdx3E2rCrspO18SSURqIBqN
ugVPp7xr7IM4RDUNv9bJ2vW69dTkDTF1bv4GJZVoW0NuWzl/oEs+ufzCLZxrtTPc03qSnKZ5TviF
aty5oMbtJd0taDq2mRTXUgWQDERGgt5QFJYPxpUT07mGi4GyzsTPOoUPiP5g7naoo8Dwk5aGpCH+
ogVqHYxie0QJr1NHn2QXs9Uz3frDaSt6Spoa/zd9tmd4AC4i5JMs0aKmrMbduEDCO81mhBcMFGkT
d/1yvU+FWo3xSEjhaGmee8FqznkY623W2YReHzLEOmRA/8KsPKbGDWdeM8GIIZJ0y0vmwH/GsgOM
Aq66JIM2x3OBgG3g4jz4uEE7LfyyxlG52ACF55Eg0oHI81amL5W2ilNWMYilXZBGvXgpSFLMSx+n
/OeCatJLHNvR+++g5HKRbpFSEBpflL95pjdHA4SlrvvkMaoZ0bNLdlcSPwB1PAXRQlBEPrQXz5jw
kOOXAxWYEx3FDgardU77CNKnPseUEYkNg3WBk90P6EHWlz3t9leb6B31QAxABLSghA96+U40o40K
3HnSS7ZdRgXH3yo6ncMNtI+UzkMwh7iqKGXFLTaVg1P7SJ+qmwGSH42QPR3ufkTtiXjsrUqwWTtg
tFduVUphObRQHTAn/J7HOu2BMEkk+Br9EHlqcI8/K3xwCtxoclxFEb8BNovWw0d3VHy1qiafVTx0
4EBz1Fsw5JFw2dvfVqUMI0Nc6/tUKjYD71DrkrAxhTKbD9Qebbu0vDOhJq+37e/rKh6WKI6C9Q2X
AGJ+hy5I7rS7WCUR0ycM8I184LTSycGhTI4inyISZu5W9Wpyue+fqOjpPMIAns5hVCfQsfC7KHYy
g1iFvKrLpwllMXxdz7o7lWlAt/aOjroJEFowzAV9NNSeliCWiPhQR1iKNIlODr8xDHAWz3RtumiW
o0dCMNJZ2LySsRlEWrYNVbE24cu6Mjz0fOkCQ67sLG14x5LTBfkpiON9DoykioC0Rqm8lOPgmrZm
ZHt+MRZUskX6KvsZxELkmIxKXBBMp8kUrrRSrF1WoTgaLRs07cvZF6D8I0C7z2f3R0aF/ViY3l1+
ZxaOpVNTwOnz8+Sf5pRmgdqR195CJAufOR3g8C3BHsyNQrOTBEA5Z/innnvnFfb3evUL3o0IPiAB
9qu98fC07MN76hWNTaxti8Si4yYs30KDkFK7rvj1FcA7MhDZzNkTJmpHe2+C6bhRgy9XHm/hhRkZ
VgHsP2Bn9595JdL9utC6jIBF24/X8JGPzxlWvc7uCCJjEJMTdiGWgjlrIR98ZDjL63JNz+Vztusg
1LDgDKo83pr4biunRLPTnvEe4raRkpTa6aqyr9gPGh3kVW4kOoi4wDDvmIiO02OGboQhbFpdWwDU
Q1ehGosrP1UiG6CYdq0uAa7EEZF2gjL5Sl2XsZmsz4LQkX8jhDkL+eUb4LDYjADMdqUm69+94QiA
EvmhMWNoUgWDYqXO1GCd6n3v+scNyNn/6ts6wFNKuceRjrSuuASbUxGq/s/uRTNEaL/po6DsecHr
aVOTbs493mx8/72gIMMVFvCqnGQnkTk9+9Jh+FyKkJYw4pA3WiaecZ20AAjYhqFNEo+Q5ZrYMs50
LNopYuF+VdjxMGG/3OuOkJSxkswJCh7EuOKuvi2xd6yCbLDBnKFDuop0O/6yK9Q8poHfG4XyAD8S
0cfST0nK12Y3c0Kq0f93AIyE3sRYboRmIhVxYPCYaPlKRk5HyQWzBM8Qr0MKEkoRhQShsVFQUV+H
tKAgXhrBbXOA5FgLcnYDdszjMpiliazCwZIjI6lqnFfbh/GIDf4YkiTWx+YsL0J0I4zIEXJoUQEX
PXj174FyPL8LLtGorUZvk++M2mELVQvokhozdMvp9fxtovqbCeoXLA/+1H/uJGhwQzcb9Mp1cS/D
ywdh1xl9UZHhQhGSDTbBjc+i7RPKahDw2OWM+xw3Fsl6KRCni7tRxX3xKcx71gDEGov3deIQmYPQ
vlSSEJeQGkuDoQpT7zF9iGPctw6JpTb2OHDtSNFlIoBIDPL4e4zW+z22hzEaIgtHTs0wuv307e5u
S1HsdCqZ8C1m8TR3Uqh87kMwZhc6+Bm8TAn6DGcCzhJglX+JomtkDpEU4C1H6m+OMsqbPRDkFV0L
3AxH29CupfyK7UEUDiIhgJmgaaDRueuZTmiJT16txd2dRTsvD6MlMF8yjuSAefcVsc5DRD0/RMYE
CAV6OaSWtpnz8ggvrSkhCbp8tajm9XWzMhdj4S6FTzwHvN0vj7TufUt2QvzhoPIdqjnGeye1/E53
yN+Nj21zVFFi6wx+zr0OnHBYCCuH39u78GG6tG68wxiG5rZGZlNXULtsjn4ZnAN4RTfW+GJIfJLa
KG+luUmUg2DGi7EoANuYAcPVoGjHCWQw1cSQK3WQzkc4W8gLOfu72hvWliENZpBy6TsG2J+8/dlg
3Xr+oj22Nd5kj2+DLhv2SnH8EtGZFMGN2TThiQO0EBF6tqgU/3LEcJEuApa7MJu0xrpc5fUHvyhz
OoJTjDWQseulYOUty+LdiEvRt8ezF/Jtx+px58Mw0xC6gj2/1OEButPruPCgbp4D7ORRcW72SPk3
USePGyKtQhYUJ3HePbzEgPHUFyewmqaW94Lf80lFXOhdaJCNKIhuLCO3y47xFVWz+KU+TWDNlb0Z
v7VoIyGm05kAaFOhHZK6cVRRIcEubpg1T50qWpI+o0tZu5ljewUd9QVtw24ypF5/bNl2NtybHYyT
XkktC9TDsk/hTNwzseBwXNItL5C7XqfiDhJpuMflOis4WnWCkwPlsAM37+xew1IrLNlwUb0RexKE
feTqXxEr3ZJz5gZ72zBXuf6RfBSxzBOHC9pzWZgb5FkrmDIxdLZgSPORlURdWCAsUt+EHsijV6GE
+IaA/TzjvTV+TZG4X6cj8ZzshX/Bh0q9UHEPyxOlX025r3k9XWKGKjp9v24sfimwHl5Hf3v0pWYP
T058ALzuHScpruLOaOM4zPePvM55tS/6DIb7Iq8crKSZacH/90J6G/GinjTDMqtlGf57d0xkB9qu
R42t2VFbwAVKEiqDLx3TkopdTY5ZBi/m4TOL+BBzGeN8gmFi+algg2IeAcS782iUstemHIXJWX4f
+DlNneGHqmERQ9ve++uovReOTYyj+OPZawy5IDHnlNEAITLEG43YtKEd5U6/+me8zl9HDYWLy149
2jy1hpz5ryEm2oczYDd4rfXh8Eamjits10HuFuzTzCoXJnkf+NQu9zY9qcXm4MBeKrTcoaNPmgRS
d1VmsxTy5qioDDVrm2OzeGpJZVRhV7lWE0BXbH3C7T1C9ehV+2rHWZhkeRzD1hEBAu6h+rAn+McZ
PTEZVeREO9SH+cjIPSZlZ5h61eibMgmrnouA813fXJMmcM/r3rtIYUnoJ8XwaxvoInqG0/GY71qO
4SHNTOH0LQtCCgIzwdtREYrLeYSpV9ZXslqm+R2znCd2ruEuCZJ6XLdVgyi9wahb9CCASAThslBJ
hxAko3/gs1omyqjAeE/FLvvIGYGtxV06/01ZYKeHJgapEOTKzAoTZ7uf0OArajURR/UOO8ma4DXV
3aJncCgwh8G4rGcgBAcHOcKZeo08pimz4RYqV2SU2SJd1BKNLraAVVhGhRzDAARNLO1BsfMiDOia
4etRWb12ZbgYwTJAs5TVw0NiUYRkkRUMlNMXbKuzs/dHuBKl/+XuGO/qILdw9Xj1RKgLJUoKw888
3u7/KySb2QSe+F2NeILiXsvzLNKWYJxVhBf0Ezz4s/79PcodRTO+l7th2jai7W6ehEVJT86S/jZk
92YRkIx+BSJrsYCplJv3vleTp9LS2k6/VaWzdQZ9CoLz2SWBtmCA8J+EZs+eHE5aEeypy0qcMdxh
xQqumd7obFtY5LDA+Jk6cricTVbEnNj5nJ7iQpUqHHCLhGX4q9eCKt9R8I97OAjEBaSsBgoZAWR8
n1aSuyVwopLGJJxZwrZhlPZj7dPzHMg82+J+0pZA/hcL062/5Qk++Ox4cWG2qthUbfA8p+vuZkaC
pz+pzvBuPNekkXB2l47H/iREAlY1493aBwI6cbOh9kPk73fJ2/+/OtiNzUfCW58Pfg3KvvtMcvVr
5tWtL4We3KD3cw49uQr7xgxELmwtgrT1s8wzx0qLIGTOftHmNYmTrXeZCxPcE0IQtM4J0BFAggWH
KHisGPUsASqF9ZnR8Ad7KNa/ZDsltgR7ImjtOm/5yPD99QmXxMGvnPYC7PYJdWiYMjJlcqt3NaU0
kNsEKZFm4m0Um1053G9MoGlwwX/vCZ2hmnbHno3Bk3uBYmf+R+pHrzN7UKf1LLKVcnn0L4Qr7FJW
sV48y2FGwkZZuv7D/cCrh296iD3mmofQa7T5tlZAZ2uNvVD3uEKx/jx5n0KYhXBi1udEVTH3DfnB
7dmKp4DzoKsYAKDVLlZW/fzIa2oDqHjChKxUokePfr4dA8FhOt4uunCR5kmdLyutRqAb+4Zkgmwj
3iCYNuVUqLiHARd/bbSTjbdQpSM54u8Ni/YkYcT5EMKpJj1HX0QXEK9889f08uWGN1dAa1XgPRe3
0HuH1EpRNOhpmHaDRuTcrvJiWE+5IBlUfSlN+KXx0aPRMqMe+E6cRSv3sHyjt6o5/Z9lZ8rhAbFB
sz25GYR6n9AfGmdMk/bbORIHpwAO6vugc3BeF03TjaV/xnG2OMuVEAdedip6vU4u9PS/ZH4ugoVl
hHslRa+GN9mqFs0n2Nhi/9IlrwGFksNrAU7m6bjloOacMfVkP86u3hpCFJTU9Oni0oeGpv9RR60T
oVpgHvB2/S7S8tJNUZQMEeW+ncEPJnNNWQXaZI19hw3yQbTdMyyIFREy3NnyIoYgfAbI2MbHIo1x
kz8a0pBNBJJWE8gC+o6PKpQP+CNNZcKnkk8Kg3aEqztgt/BXtAkSU4kkEhY1Feh1PFvWAepstrWW
N7CnzRshFufvwn4DglZbdaM0bpRF2d7WYw2R9uBQaCuWatUV7xyjLSqVpa/8SiBIRyYVXG+kHTUg
o+1229jx+0KTyk0+GZJnolo3bejq1HhgmWTYJxIBwlYValXZDpeJVqj6wR6m/G32H1hK6ubi4gxp
iBT8PzXh/xYwUR4e/9d9oSYLtDvatly8LSo+fgIbQGy6I2PLCTlREz/l4Q2YXYRWe5CQL8YAZGnu
z1xveAMvJ2h9azFvETP+zJzB9PhxbGwDca/Z02MI4VLt1qC54CgpNVpjKtnf7lJT8HjZyU2YT/5w
dZm3rYls5myW/xaNYS9h2YA14pWTVN7cd4sagCbtiujDVBDPFtjiF//SdZT6EEMX/HT80YGXKkQC
dNRdwW4PQkb85/beorVIaRIbCl5LNgecq2Ho98RdQ8ZhrMQtJPzXicI0NX/r0hKVOM8a4WjimnkE
amu5KxSmjbDA3vro4lSknrl4ebyi9qj1A/X1zFiTKhWG5qFUkVnW3VjUkTjnYjvrSDUT3P/6LVs2
DhAZ2A0m7OkjFxTryojARzYK50IoCTmLNsCxstyUVYizB1RtIZoF+Qe3UOqYtmy/kftKkwYxnPuT
wLfDVFugHAFn0ZOkUl5sYWFVXn30y/HEi2hbTNL8HTlTt34nJot81aMjVrrnqYQS1aYATADYrnGd
ZJ9UqLFIxuIbX+947qzLL3tU6lhVjFdQtF+PwM3sENVLsOgLk3IhYe8bLEdcBmO7etNE0CFsQBcE
6i0ZgCXPJBS58MdW1/ps75nmzjpqXukfvpc2d5v873MsNhgNIZgSHf6cWgUXSSjpMqu6y9Ksc7Yb
0s97i8wI44uQZSHxn1gfTNgi4L0oh2plzQDhFVriwexSDoJXW2VRvojucZWdDR+fHB8ibP6pR0an
/BE1pcfzaHMXzjEMGxAbNu8CIEN9XAXruzx2T2mvS9DvPcXxYYzDnWvsIWuVDPRjx+p6lZlmWZTC
hhAnnl0ySer2S+E9d5bTlsJvAYC2/kt58hxgRYWMO2jeP/f2I7j6upJbsy5U3tfBbRbg3DsMAR5X
D8KgQpjLJO8iyPV4SS6FAwnQIwwWYjybLnpGih+jXcV/FAFz1/vDizOwG7z22qPv1c/G1jZUBdgy
fsUiuwuXGFGoYciHbGt6kQ9vH6M+hArhh20lTetWwXfT2HqDM3IIyKd71WZpS2G51nC0E+QLFIm1
Eze1vV85zVi3qOlCZ9Bj5UQvdD/D3roJvJhA4lrx0UmS5BqTqBEiybWdREE5yrcnb/s9Vgia8Bp4
pEsTZ7SwuGH6ZtwSzjXfrC/dOwXKCiZyZ1g1UP1JBugmVd/junbCa+rI5JnWF+pJtHDi8UVO+q+p
jF6FroY/99sdPvoN7FYnRJhrQxe8o8xyoI5pDbWUuz2Gw1ABjJQSoM1Enri34xjuD9qtsilSda1c
9Jaew5ZMBe1EhmlGKtl5VA1y7LjLnaHOj8QOjiFxlGsqadL/EJgMYMjLtNnAKgxSoSxIuJ9yvWgC
QORBHRF+DUj3/LZsy3V3myqPkEdI0KPGWlAKMl0MRT/AHxdp9FMeMFJvYN0VIhs20nqIZFLq59PL
SvBtW9TeKgayQIo9hECvYA1abcsm78MvzJK1ERBCKYNqcaGAqpvWty152uP87k+8ro7yv1GzReh2
Ryo02KTZQR0YcSc4TvGqYTsmNtDN1s3NDb7a2S0dAY067gmntDkcGtH+iJ/vqJCrie8k2qwPHf3S
jwC5CGXM5Gc3aLSxfBjN3EODVKoTvXOiiH/rhvW2DcJ2MkxAlp+ECNLWdhOX87pz4tgmM6tfjAXI
wHZo/bOqD+soFvNwXN0f5Qbwu3gz5EDJPxNeXgl+nIz1v3skyrmOWo6yJU1vyBHA49MWDOsX4dqY
OOwCB67DY4rn46BUlboWHtpru0jrKD8pKcUh2prnsqlD3Nf6mXJU/D3Y6OIV+/pFv8+mz1OHRi5u
3g1KjCl/pIAFmNDolZ5fESerE1MdrJ33tVRuB3ZzHvpX93W6+fpG2X4+SalOxH8ceL3YOjErIinT
qyFxJUbUXcUUuqdnHf8Rs15nW2RTvMOvep6+8lkaHhuHCRYb04UIBhc04dbr5P/97S9ui9OJcU7u
XjIE0XqyJVlUUhcnlszuVQx2B5L/dhe7IU/SX0d6YYanAPoQFXANJpnWe0j15JNzIeYe2k9EWXdB
ZU0ctf8F/6GvcNQRcGBNknpbmSyG4E2sqZ1mGOy3DbrqLrkIwWocYM42nAjRh+3IP8UwnqZUgm4M
3uPK8Db/KJXqTzswN4jgS/O4smxI8iuo2PDA2K9VBAveCN1mE8xXChssO9dWYk2OUfHoyn0OZ5F0
OxtWAkw0Dr+YXrGjkd9Ffqzwfwc7LlMAfP9iwLVjldiJSRwujIcXWy6EOKsHhE0y1BDMoYdyl74H
4w4zuBHO9ZR1oz+M+ra4hC+QtV+TW9ITuY4zWOeQdj3xJybRK9PStEKpiLIr6jWDXKAvb8Mcsd6Y
/elX2aZcWRnZknMpa1qbKPkEhyJxQfvec0rZVqqd+2eQUCeTwahINv95JTyfL8k+lhPTrS/a/Ts8
e8fmGr/brJO7oFPkUbtr7fYW0geEXd6kJxamdnwaF387KZf75LhT2HJXo8r3iowh+TulU8tmGApJ
k0gryhrehO+Zplv7YMuwWSlXAv4vKfUvWIfizittaEKR2bHIQxUXC0+OPbo1DN9sf7FdzPqYrY2f
3W+xhjqJHzWi+ybhfspNidofk51lvRQQstBUabW8zz9H8lLhY+380dK9irqJ989CVwkh8+a5Nnx0
aQiAVxGez7NqE4Od76dl2BmBuJvFW5057kf/ndEuzgnSFiuCR4R/D1Cip2NHgYn/qCnlFuV84UeJ
0NoOpQnpVQZjP9Z7CMtTSuhd2mYnDqOI9M2Q0qbVRl8lVbBHoypOurlLkUEWNmeI9Sn3XPm3FXov
xCW9l7XALwYZYTMkFa+u5Qru6ZyPnrRrw2JjUtPjFNKePKsciC7qTYQglm1F7vaasG6simjYhoxS
ihXVpPDcd55uduoxWGrkyr5POueDupIb10HqQjx2zIHENZXTrMAg6C4w2kcyQsrntTbL+jqK94d2
uveDbbjmZW5pT4iAqxrv8pvuHJWr8tz7OpcKKXqCWrulgwrcAg/hEHvznmpvAwuYcRGCogFGGVIr
E6EfaT02GhOo52DZouTWmEgGg6E7wb/IDQRSkdWAPrFuWDNzpdaSdLueSyUKRjF9p4HHVjg8mMkz
sK0On1OXsWrrwP5iPdv00wJM8aWPObDFYkcmzxfoNTAFYAIsUMgJJJ8rpaUZ+Fxnwz18n7CpsNQ8
KQMSouIOQ6Fr+1eghnQHn6OsASIBPI7rheQwt1saEb2S7z+itJapztnpLeNFisUUy5G8wOQhxi2u
YsatejRBa/Ck7svLrCdmf/6tsegse5EQWdgwuVTssV+/P/JckmdDcIYpxLKbwfFSAjnzogxib1Lw
D/fIBGiHY2YF5sN9N4TCRb5bymx4b/+avZe07y5NNhtMvKaDS3NhyjoEYcxqHMUiv+tcs+L8kEny
njXquxsPvHOx4XKyFHn6ucnr7MRIKdOaKpq/2IgSXJHSVOgKZ1X07Y8u/7mC77GcrbCZX49dBfqL
Qnw1SPXEfIamw4LddRPVnJTtAUxZhO6+Hx9oASuEjUVsa9SOY+Mb7Usm0zenc6cvWApHdeH3550C
m2hiK1ZOtMWZBNR4VF1cN7t0Ew7Zf2YeOM/5DdfynpoXxEM1MEWHJSMR7IR50pwWuDb2M/n+YMgI
xdez+BRHk6JKfQVr+sMsTt0wmNBEgQnVRlVRbguRMqFYpcunJ2n0RiFi0mURnBLcQioSomGXPLVn
oXxl6S8NhX+sYu+BVCfq8CFbttYhzPsznhnfEj47VXFX2FlVKJHhOh6kPO+7icMSyjpgHJfQvJub
BZVOT+hMUsb6ktOktI2gWvl5RzPRgso89+5srfSoNxTL6rFqr0/6x40uKitxnNam4Y5bEA/fq100
T2eapTQEsf9gcaozcAq4JFv5tyZQq2dc/WdDnf1/+DlyDs+jEqLJgBX+/C0SOo+lnp6gJ7nigcPe
BkvA6djwchsiUGS3M5z0rizx825msi3jgTaEctymO4yc2fJxdCxrB2IUjgHlU8TEd60OfU9m2iON
zKkS3KxUd8kGFCHuapfAKJlMGdRVddRY7VO7QsZflcc+ZPfdZ4zktcgxoT4YjGZ862xDGHPUWqZz
TtQYGAl3U2sIDIdZhbqOu2u6d2LqyDpk5pPUnEOZkzskCKE95ZMi3addzYdggj7CLi9Oo2tnf/Sg
AcZ3yUzAZpj231kNQQ1gEPvZnbBBCWfg3zO+RSKXV+VJYyz1WwTuH30EBid5eDhDGiZnIIDFJG4Z
cCoeSRBDhJRppgXxB2d3YJWi5VFPu/0HgbvvhQlZhwPVhcjUpLhyww1UIbDcK10wEkicawskvlRf
jpu9IHM9GufkUewZjO/HRqeQhIDUVO8ZYdnpOgJtLblmDrfpOsPuVyZUKXlOkpsp35ryII5hdxMs
BQ/kclS+UCqfDmD1m3G/APxglbS9OeFLr/ehA/CSx3Azt91EyFmN1qM1u6eC3E0+CRxbzx9srk0i
q+NyQV0NDl7SdUo4Ww74vfMynRZD2h0hwJ7xnA7auSmqqdnhUMy7aprLVAJYSH+IkeWpub1Q738M
xgYmLbUu8Wnrf4HmfpFn3T6ndoRUg6l0T3Xs9kkhfyaZdgCZsmoYOoqC4Clqdp5UE8qeOG5oxKFz
Ee0bdRdijHAnHWsbPFEJRf2hQRnTmRE78b2/sovNPiVWKJlTteLQTFon1vvJmhPBT/PaRNoVItqa
DD1fpeiSyft7XK9r3hfc2TTl4UvUmMQYX2rcMYP4PNT0+UfGxvL54SrNao63RHELTJmItccwpjZd
yrDfWRT3AvGbbmFc4DjyLB99YBxKLbIXZOuqK0zkYDNsRj3eyPtr1SxewjtVrllkOzRzrAjN6WCg
rRk8GMmNvDYWhArfoJAfi3jywE9u0s87xqhnzFt7Ipm6/h0A5Fh3pc751Yv92IxSz+Yh0DVbOWy+
cfWtjNTelgB8SKiRDmiRcWu54KbwKRWjaTy1l5BW9PVvFw5OLjzFzraWehPQN+NH30IpBXcF34Hl
unq84y63d0Uoni9eF39a9o9hhSh0cYi7xm/O6tdpBiRH4NoQly0/Ts/hlN4GQbHphEnSCa7WM+yR
9TJyLPjH14gnGST2DBKanGjtbTCdLlJNq6/OWQoMkZ/qOAYxiGpg90UTexvvVoyzJdnDC55ml6oJ
EiavO5tNwl8IReyY20kkymVzK7yUwW5kqDEFe2nMxQBMD2drgbXN0QEPHxodAyOXwQq5cjkgom75
5Q/8CBEKQHt3T0EYKlNeAv2w+WMelmyhiNnujmxeHr6sogJbGt72KxXAs/0qLgdbzNjdrCcTUj0h
uwaEpix1TmYw5/VMGzhOLcK8cClWDe/kTmHSxBo0spqyhDjAkBb5D7vXoVHt0VzK0qzaTEV+iKeI
IrQjwTeQf45FW1obw8Mr+2rGK/lhgGjYb+6KAVU0DswrjY5Pqyn9G8nBePltK/qJHhxVDX2MeY65
7fZMVUotdRGNgBFl4zXU4ZBBXSXe5SZVVC20F/leHBuBngNWTOZeYUhHz3dHMmIz7Yjo0cQteUBt
wFleg4LeOyY9GLGsSHs3D0hrIQkpihGBR8LiIDYm5iE0xRgAH2GFmfXvE/+aqGyZvrxecMm30lrS
tvds/DlWOojP3GAgiSzxH9lV4ofPnMyvHV58x/LJYaN1oZSzrY0880OibzY7Q9+d5+Lj2do/HNwU
hjBdE8d7QO/69vQ08nw10YeLmFO7fW+yxBbBJC2XbT1BWMDO207cguqDvpVELvaEXB5ZuywhyW8k
eWksTRmN14KRss1dMg8aakKqR//LBVIlHGre8BReJtW2H0wBFDwuj4q5RZLmeyOgtgV3j2YIIuwl
Q0AJ5azcy7847VcFqqvERMt9zzxI/DNuf3e43hYP2+CfDKixn1a8rR+knY1pBwmCgdvr0G436npQ
Fyw+uWWKLQ/1mu7mPeg6IuOncfuvyDOklp5lf7KpzJQ3kjTSIwmk0RGI+dTYpC0LpmhuN2F0KrEi
LHkDjn6V+q3yRkoX2FGQCyd9ZUhiFMRGhbnBQHgXfK2YrE6gcvmP5O2Kq052VRy61I2XC4Gf2OCH
DigCymMaNBKaUBlObMXE/9dRdo+/EvEIVE2Bm0iMJcL0x2Fvya+YzRxVcgvsZ50VnLLQGMJ9ZlKv
vdJJq1Ko6VPdFoQjUJkgj2+Tbnp/PN4upfgn40PXPc1XSgC3Uxo1vy+l2SG7KH6WN7ZUvZplMr+Y
/toxOSXqEGlnFhDO6mbPwmwoxKU/6BtAOcf1dOgEG8IBladlVTikKZxDFxnK/JdFWIE1p0+0gpwj
iG8GvI7PJVfFz21afyHrtW/dVfRdX2R9T9TbT7HG3R5Pue19fm3PRncWN8jBSJ6y0PSx1fphk3ly
DhPqiWdmoxW8W5jl/taladSCVthYeI//INcx7RwgomPQ+oCW0rFpPJfPi7l7R2DJnT2V1WckjGJk
lxjmDDpUP5b32kW280RmO73X9Fp5qPKtO06rQXxW2QXCZoRGNQ2y46mvfTsGQPKdbRya9aM8yvj+
kKIpSrUEdFPTAhzAId1He53M3HpgKpIqIcSVDsO1jT/8BShwjShqhnhFBTZ52wFeQY3vNWzABHgJ
3gx6Q+Df7bb2q+vRhTs8NYqEk5j0bk5mFoJjh4ZUvL8XKn1vMJbnHIxf2LRx6OB4I6g18pdOrbwC
Xq6nkmNq96x3r5bV3EGeA2KjYUL5sNywrvWKhqa529hW2jSp1OS5/uPk7VHqNMT+R+CpBbE2P10t
pRqnuNxVtz/N6qz/Fqj5mQeeL4t3p4r6bUfHLQ5NHmjnPzPo3x6W/Lz4bil8jDQRqOTGjq6bWSiB
c8/bKN/XkaQWGoOQIxIeOn1rVxyq1CXYSR/p7y6DzMlrQOfyNM7xYjnGVBc109tN2u+2Xse/nOes
34GUlsm3BylqdznA113RhDL6u/sJ7mWm2LWzYYdA0xoG2T54uKUGkPJ59Vskr5LKU/6FspGz1llR
dTmU+4Hc1+RjaYoy4UCUg77+7TRwlrbtQgc7VPEhuZvvEN//Bg6yRcI9cEIJ0I6+aES7jXVmc1e0
H0R2brYtYyiqAEBQZUjtT9v4g6E9QkzPIiiYLTKkc7rcWbXou4ntM1THOm7pTii/3M8bVLzMyGge
oTzZhc1fl/uNy848G70roVZQCznOQ+VIGZ+RzrxL1IQWkwy9e0HUmGAIRi3Ad7lXyHoaDX4S0ftf
WqSEPgY284jC9wJ+c6PbggUqh2ADnf1o3ntsryZOcJIt0qdNOa7xurxpN0fs7V6Cz5/vveXIRTbz
5qLcI6FKKiuW4H9OWbqbeAFMLnDWIXs0VL9DDjn2vmE+GVcRZUXWmqldZRoIzOjgMTf5n/fyoPNL
eWgZD8Xf1D3yww26ueQtY9YxP8utXSNkHcHQpc/4EtUEyvKBRbpl6fLwSna4mXBkYvbCdzClHroW
gcCMyJ9o9pNq8xvlJOdJxa+aC/8QK35DbnDsuf6Np3krwb42XXdFvVz3Tlm72FtnlUa8iGCmZmtJ
tX+5+u1ONbDeC+WGa4EhNAbtl3hev1nhGhvk68qJzA2hWDuFJVyWtJaEQ3jQG6kzrNtyppKywd+b
d1A6TXTDMSQ7vpCI5rc/6GqrrqHuR96wnx0MNZvGUTK3wksoD6QCVuEIrmMqkzJY97MGcgksDB3Z
O16tDCSfRRjNelFFofO0jAsRMJomML4Va5qi5c7Qb+9Ra3+/js8BYvMFAqt42bjhk1+JplW6mxGx
39w6Z0dTyJDNLab6HgVCE1HFg5VaeD+vhoB+S82OPlSzRCOT4rQt0VTgbdWuLZIdZtp9mTWFNHJO
euNycPOwmzY/9MlJUUcPKmYOUwLWh4FmGkOIP7pJC9c/4XOK4PP1wSzI2xNk1QXHHvC5l/LBjala
nvxxlq8WIxyLCbKLmOPpsKdCLZfJWjOYFfmSfbTAbQzjZyiumXMT0q4sNkjLEfdmh+lD/0hYRmCw
j+EHwC9d9TELopHd7TasRcyl1BcMB8adIiodYNL4BwfUnfBHjCFgmRZqcJYgI16rAcI8n93bAVkZ
mzm3qEgNK4tMHIYyi8GLHQH5y9pN2JmxJsvmeWPI9m0QtwnmuowyuA15Guw+ZOOiOF4sAAo992Fu
owTDhHWqKCVJlRKjWGDgd43xvw17uk4JQ0aJjl2cUQSkDaH3Ah1Xsfwgv837WtvylUShwu2DUhmh
0JRLHIEu66yXam9HNcPEeidrlZXejEgss8QYp0XPLBmCJpr4VHm8soPiHeeddU4C+10sz/mabncX
Mzo2lsgEAAJ1N6n93JJuDmodyBdQCS6bIBuAN30c1rSxjQex2r+lOhfDHzUmuMzu7ZSGxq3XGyS3
mw+mKO+h7C0eOOViKpsgeql32s4Ufm+qmWg2iPh3ldqoet4bakHzPjhUMPsPoie07hxbS5YzCwd+
gU0kEr4YGgnjGQSUiKIoIRl43D4QnAbiqplg4WmDxoe2/qR2h3QGG45lW9Ql7X0Mca9MnKcP4Qof
sIgurXRj024s2g6TxlA66XOiDdu6blpxhnzGlqp+unlbHyV/HkM0yl3fpOlVByJkEVMGPpoI9ZUz
OvTXCVxwJs85aF4IQVywXAZFpiU4TwfhEWIwsj6vFc7mv9qrP6qxeoTUl1eVJDRswXYnytvUyI3J
fiiQBt9Xuo/ppBBiPxLn5NjlLYXhpHogKcx5wbYJFd7ZRtQb3PDNpScPKPbXD0qjpvjRtWbOaagh
Ac1PcEkmyFa5eSS8ZyNYc/MOpEF29tT+0JEUdtJvkD9OVvqm8+eiAKyL659P4BUQ6J9CbiAQtY3h
WUxBNu3Ppt3okDtqBM/HaU8KqLDiVsryAP1F5Gu53t+m4S0cBK8Bi1Adkdx2lIfZkYY0jPvsF+W6
gdrCah2lBwTxEFpD2+/MPQDGO2xSSLvm2KiQXZQj8FioQPT4i93XmivRP6RYP4Zp4eH1KtUKxoOI
QEzVZPkhBweTWLGfZKucmx+4dzbE9y8hYbDy8EqjyAKR4Rooe+icmBhn+NCsjfjc5qvI4ZaMZGK7
G3FBMRxlquk5FtfWsDwICp5L5BUHL9jduIzXBIn1K2vGsdZlcLjOVmaB8g3mBPVQ6NkPiJLprK9W
eQtjxLhKjY7LfiuyroJBUO486Re/+1KziZp5SQ9hWIO7jZ65ddW9kQnqAWWfEeTNcpzb67lKK8P7
WqvnZ3cZyJAsUxuaWqbZb7hZ6d8JP1vx/5bIZERvpnYLyuRkXsWtic4Hul8TAytoeu2YBye1xIgp
Bb/VteSlpPPeFwNhkfwNBjnwV4VazX3ng7aNrwLKheY8uQz3buAFGjNNHIS2OVNUx1QyjfknGyol
WfcHfhGzXGuKCIl6Ckr7gylgNLhzoIEVFKPiaF5yH7396QCAcE6I9wD8xr3DxQK6H+0JNeiIa8YU
H0+I2l2BP+2S2XIrhUJ6zzkyfo6w7TV1Nb4MBC7fuC0fqP9eQ+v8BKLgbaz7TkAzShv1qeCjrqAt
hcYIvX0sLiEpSWVAftw6Z94YTSIKO8b3xFP2mMQmBiZwRajqgx7F5UI+ynWMaFOINdTb7MOvIAwi
C2S/ySsi4VQqmvja/IfvFsV51Y2YT14s4LYLhcwR9hzNSjGQZ9iCUN+WlxPDwfmRzdEnKwN/BxY8
YEW7V1y0eeCjCn/g7aS3wXLbRWPzhYEE9fxJXsI2vdk9WsVlOToWAePLUr/aLMqe0IdJfXgVEzkR
bt/O5YXQwAC5hz8x63jAGj1s9UnCZY3AyEc3g4wSUurT8xIoeCn9Am2otsPrX4sNbsChXDHzTwxO
UyKdV1RigqP1k5PK84b2XgvMoTeLl/z42FRCtybwM0qs8w/hf8bZw9ZYtRQ03objROy2ogUkncng
cwMocybs9UGL8xro0vlWjNqrZM6yADg5yEcm7xwNJLuXODXqbhBocf4Higk0fooar1xMc/OXMm13
Rv3lxztpyS+Vfv+rxVIS8rdwmkLLgQiT+EJzTWfEbXppU3HgL/bXTlEO7z6619pUWl/ezf4A4gBB
ReiwYX9qUvX8iYA3pHaT3qRuQEBrhl7+KHBIK0i/CaimqA7hggBc2sdbPo+MfLjonn957Dpf1s2p
+TPCSC2WOaA0XjXbcacFe568/pGaBEuCmyDHdGcU2rNvIqMHeXTuIQzlUJtQp7CWlsRSjpwPwpOm
0w+3pDsAaKD4CVsM95v/uwPEln8/pSYeem2cUGWsxCMwEhKMG3ayPTk/AcZDPfzgJNiB0uoXkKub
Zi3nI1nxRvquAJwPMDKZSra3bHhxYZizW0KeQ05BiDyqI3ZdzdPqthoLJZ0SclbTR6xrsV071ypj
BrfsjJT7jZqK2npqJUT3ZaEKsVr1OnHiqh8xLsfbT5HqsxkILX9nTCjvHM005X7m8HbgL6g5cqv7
ikn7cUSP8K3+22qFDZ5AZv9VDmncSeUQwpZJOWVWdWBIFDOX7FB2Du7v5DQaVtpDtUGhAynu9upE
EGZVH2Imo2Cv8BzRJYKnR+mNxtZARd/GLWTViXiP/llZdwcct2s7/DF/140G1bXnH01cGtiH8l3p
Qlrrd/YKSqwyGVFwOLarxmHyEM9yW/HekqqGKDt+wRPcDSQRwgklFTlWffGUQ7iUQLu6TWU5edeO
7aXuImoaymN6bWgohAvQV9eQS4w0G6yO9w1aLr/dCtjVjrLpXDiR3/cEmWz7/pxDrpMA0IlO935b
j2b93Zs2CvZMley+BYYmZFHrHr2tlMXNQZwdbydUJWge9UvYHq7aNHPLi2IzAQUXAOhLJ3fc5qzh
CfLPCpA0aiVUsumuc/+vDDejyp9ZsgJ0PA043DetqPPO96GcQd5szQTRiRaEl1EWignC9OMgIO+f
lDbFBSqsYRxAnPRoWS6RfGc7z1R86pJRpwUN24wnjHWvCsqO9Pjxb2SdCtrHiS/BRu1sH3uVG0tn
dDA7mOLpvURtKi53mj/oY8YcBbUmjqpK7ZylXIyXLQdVt2bkYLMp2cQepA==
`protect end_protected
