`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
k1TNL46COhbmajA5SKRiGL/yY/l+mDLK/tFf+4A3HrKrF54pGquF9pt8iogqr6NpcWrTvB/+5+em
uF3qey4pJA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OcMMrdACL1+XI9+3IL77pujXvR340n8QPsMSnO/2DpRK4Y9zF/C2zMEaC+5uxqsE6PwKLSXPzeF/
IC1kWxHQKxI5mk2ZeBSsrFRL5K9uiEjOODHu7ANYk0PEpzAPBj1oKaATyTeE1h2WCQ+08zWbU4+4
//x5NvPGnOmpf3Muz54=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
yV1s5CuLMOTxnsxqCKPOQeVbUNk8NcuwNdhjTikrBhAkcDuYIGXojoKVM+imIaAyGHiEACHH6Ps7
oi+WoWuplClfWkapYIy28TfkKVI83ukfoc02JKrT3c1GPd70i2IloCqFd4haKR3hnMiebSM4p4mV
fkcbl78dOs6wMTFZtFNIjdrHIBtoo1U9d2Cd8VkSvfGTteK2f8lZgZiLr0tbK2PDiYnEw7Pm6dAR
R7whxJbvmKup9gGUlFk8r9WhkRZEpVmmcBCP1wXsYZ9Gbq7tZidIcrjOV0id6d1IEaOCqZVL+STQ
eXP11L5W8VnodRDh58M/PDksw5YQCFpjJvl8wQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q57uFnCR7T8tBAoMNBT+XJHCC8KWAqe0YCE5G2iK8KpMAdetvYrZDijVNL79FxnPtrl0efDWj6TN
lw/4Cmnm0pJTYWzY4cdb9lpn3rbpFV0yEvHdVl2D6gninJNs0Uz2/E6Ke/cpoUfq2zjpfQ8Tzauw
WBXAcjpYo5Xiq+rsXcmsC1I9ZSkctCHZSKB5JOWh2diBmvO2ag8IncyZ8nMYSWPuYnW8ZlWNL+pC
JE/VTb1mlRKCuy5nI0rEjn+jIPjAhc25VYWaNO9nEipYkzBelLL8JSbsmBFal3yCQaSDwvSBzHbH
4aQFaK/r8V6yR7lJionPar+JhgvyK284MBy9pg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sk2HaHfm82TvnE4/afj3DwTj6+hsiujE5Ltt6Fq/jHWV2t6q59CMzsnceSUKPx4RZIbJl/Q181PQ
ZsmBTBEW9IgLjx5HbJDarOPOz2BSRZIYweKp/8AgCCdYFaAAid2Numa9hGNIMZHX6lEulq5RUE4j
Gb8/nuMc0Uox5TAAfqDaIv7UjUKzaFV/51e2xR3Q6F8Eo4V69ILEHi1N8KepggOJMF00gxvfBbBd
dRKDAPnE1caVZH9Xf42/T+TM0bAwhIfyObwZJSvlYaZceNtLmdudMus9y5jJUZ4Bop4ruUnuGTkx
6q/gbKPwmh//xaA8Hr9rOIz5Ayi+4+nGkX73sw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
p384vz9FHp7DCLW3O/lTGCxfw4G8ZO9oWer4u9Ywwbyzotl2fprbbj//scFDtINQ9aStJOveSBaD
8zx4338oQ5sqUI6+wNoupWc0RFhivVayYKuQ+eKeFDJWQ9eRzBd1iwoZh1/D5/4FzRwFZ52Y6Dx5
/L+yn7KmTMdhpkpwwPw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mvIqzEhj8NgcfeaiFxhx5YejknA/JByLRLxkd2+a+A19X9stdBHzILcp7hfD93GtrbWwYl+rINSv
qZqKWfn4Z4BqupVlmeItUtr61qOV84gMONb4FjVlbygM6fR+jXRLjYGNuQri1Jphak2TPa0MdeXP
YXJy15KUegyU0CTLm3nDHVP0YkPBAAnA2SQ1LHPZmVGYB4RJ1q15+2Awx1zTXPyefMda3Va1wlHz
GdvuKyjrHgEVDz2kSWSZei21SybMnl3IY0ZkgG6ckt+JOtyIl9XEN21FgSMA0vrP8cEwfxPC5PNi
paQ551BLPLze5uwnbrEUELnVtVSrGSD+GTiyjg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 170448)
`protect data_block
ECJVlFcwAZH7B7YXvB8HnAL0ZNFE1AzCMwQYBbF7H+8sqcVP1qHbvC7ABm87je5KFHNJaQBEUTjV
Fu7V6cFPhEBu94yoxBMJm/Xj7BESTkwA1SEavuKWfVIOU/VKCMxV7iuRF8nW/2/yizy9eBPcdTUM
R7ZyugY4DA5jdS2Y1Lu+bPvDOQub3SvEQX1XLgbi+N2RkXB1KSOpHU0f8zXCeZJR2YVw1Plu89MS
Ev+waMjp+YhHjWQ/n9+Ebvg9GnKDpgJ/WivFk5zk+KI4bnvGPoYB3qLNzZ/oiJNpiRT5DPtQcAU2
8bzaQA2GmJ1xxrd7pBZkRXEMmO71G/+E5v9BqZ7L819hYooXRV7GRB+m8eaITHCigfLFfDrLhAoR
2IrkPPt97e8i3PHHpfk5GOgPrb4NK/fFask+YEa5yjzBTQG0v11coQkSTfID/8SzxQZGL2I4AJBT
jHNkOrWBNEuDnWJIdMP/pc5WWld4WdWFRVPtnof9Y1esNXbiHHtAkoZBXS9qwN+H9QAMgqsFnsPR
xBtXRQKXRBr8dYdJP4YkHhIYCX+Z0qjGJCqzHMhMzdFYXdbBD8ChfD66fYHnk6CgSICPaLXsLdM9
bkxRbdt4FaFWZt/OHS/Gjo3EZuOPUXhRXCZUiMAJgius4gu8hwQUxt4vbCKLWrEo2dKiqAXMvAXR
fBrakPn5WA0y5ccBNX8cQPTTf+T7hZ5ysCUGDtnuRj1Y9mDUwXq2E7HE+EYv3VLSi7v9bHaL2d1G
TtUg+gdlxUDtxMXyOdT+GanX9UaKAXWw7J3RbbyJSwxqrTruGVcG7hSVW4eCz6X+swdkNZYvXTur
Rtv5UMDzFYkvxK76b1WBcgqWBFIQU3dDHGGPu0ruJyeh97c13+pSXCqKVyY6llhaQzbzI2k7Ad1p
IFbXbc6izh+0wKk8vfuwcxzfpvZsm9wi001UoEbtlfMU6lyHg6thC/iPvD3apjTCJiHHTO+PjBgP
ZXyQqhJTua9wcek//6btTa0gjrWucRRKtMyKSW2GSpN4/Edyx2he+hQxMf0Ge2RJkMBGuLDmj3Cv
AUO8iOMqqqmMbR3r/vEylOZ4z/olx09uZV6nMeR6xBVLX7l9I6kWSmZtGaHy6hDgeI1QLzIB4m0X
CCMeX7WO3lwtLsjvZOAALV0hEYt+dMJTR0+eQJ5RXzaj5bNFZ7856UZYWfjAvX/tXQA4DTNLEvIF
s2jYhhNU67c9qWgnmtQeWfF5n+nnQmuDupL7Ry1qLraZMhE7nIvXpvTRWbmAMIKtqTy3OXevbMpt
KXsvVmjxfv4k2pVjRpt4ejgFISIGL4u9YUwgR00kqMkdvGkqBFANM/B+bjvMVCQCk+YrZpzsU8s7
ZSL2aO4xldL1TqGQo5rkz/PAHI7HO0mhyoXHtzW20V+T4+UW6YP9qt9gKNfxoofUr70l8w/ImVBq
aFi8s1T1IE6L5XueVvdj1RingWo8swPFXA/c/QkrdOeTi4QU2cOHacUsutxa49qJ9wVVU/0saxzB
685UNS7WvMIV7v/5I45dIxPwIGIE4hVfbzfrX9PLyOl72EOTVPLQBx25/cmUERm4TgqMEyDQ4HzS
wmWodzrvpP2VnZrLoH+NuP0xIn9C2QuyjnIiaL3l6LtXEP6R4M/KmwdwiJaTTb/hNmksu4jiv1cw
Lk1NXTGFsxWG81kK1LWBOtAwSGwpiwzKztLI9WuMgpWVMGEgRSJfCsChCBAYHkPKSNYsTkdpKd81
zCKwd0WLqf4GQaZzgfjCP/oOTS+6WyFxca3DAW+DeH4bJnVN3nK74D0ssrrsoSRbYZU5rc2SpFhN
uHDriO4WQTussyhXofvuqGcJlsJnv2xQmaH27MXV9zI+XF6HVZCDW+9rFzC5SZLtIvQSGmGhtQ7v
6CEtrAaC7jdot0k+T8DKv+cx5uKZ7t1QBLvaRRfSOG6ZIti0VBHyn4lBhxqoWOCdwQvsLbKrzgGf
oqmaOg53dKfrsbVNYAXDgKOlVYw8k4ZkHtyrsz8b6eWAFQ7+0bIogX3aYHDqQM4niZOr5hyO4FgT
0RedOaPIHBiNySOxDStkvlR3sQTnnmHbzQ5Yn2ztXtKKQ5OCZsXFbBHjuE6D8IyKNruRafDFr7+g
eszlphMv6njXdz/O2Jgu2sqAiE29RL/dJGSuos6Ad02ugqigtkEnMDUiE/eFUdwwQ9gpyc1uEiXJ
igRsP7/bq1zDDUrRaFs8LY+o/sj7U7vC5Ku/hOSt7B0xIdsOXgz32Kvf9VSOOELKZezjyhVJ9oxv
cyyQsd7wQTmDPFYs8wKB1kWJhRONqX03w/BtRWvpCotII4OkyJMUY81gQjIYuDieZL9mrl5HLZaK
199VMNHJxDRGzy59REu8dd/Sy/QIdRiRteNauxXWRmV1Avb1IPN6szLOoJJYMtFTJL6TC8kgqt7b
1ni3wII6rcadcWyQCmfgAZ5r9zIR5I7KM+2DTWOeVGceP3H9U/L6A57gz23LCBzwworGVdo2elej
UUiDsK0LDiiwgFTgSR29fYRmvewyCZzKP8ztSoUFmBI4fFsRnJxOyl+X0V7/o1WDZYgYgciMfZkH
rSlhY9+IiMRKKNLhNxMWlHjMCFqSwHqbXkkUZoVu4VXkvnZT13ozvZTXfNKwJVWlp4A4jK9S0USe
yEuQE9JuiLeRnLBz/FdyWx0wLZFjxSQiOoErBjKqS5U38M8+29rntINe/o8ueHJbadFQP2M+fPhG
YHNCTt0JqDshwcAyJjCLMWoAbHJrC5EZddCWZoNHEjX+O12bXeOiJRyDby6W5ZPJ8epEsUBMvTba
CLZj0uqwkJmq1g1AndG3Y2OIkamQywGE/Z1aoeJMQSpoXoTHQFVKIuHJ9xZwzVTG8YObuLwv7A7V
xacBRaH6QyoKREoEWcznso1HI4Seu04V05LndXYF8Bh91kyiYsAywPh6HTarglQHIQaJMkPtWJhY
Oq/4ExunPn/de1YTuf3hFG0EL3tzTs28OXwIowAM6sGAa1IgZ2W6StIUXps1R6L8bIXTGgfi5bWo
yhGW0rsw1vmoYHVM3zV8TqizsHd0guIbTrtG6uO9VJxZvFV55+kFCqe41l4+n73rd8R45Tdx5yi2
a23cigQKYWATXX/OzTL0VLd0Aa2yhJb+SO0WyRkTGchR3aFDQp/HPwclh7fhKFiahz6XeZ9/r42P
PPxKx3mUqQY0zJ87aZFkV41T2z1knCAA2RNyQXhz+OchEhHOFP2XtAdcdTak4oVu4tfHVtIbNGVW
r76obpp/arM/N13WA+aijLXmEqchaexpzRQeocXdgHIqgZnZ8Gna8LnBHF2Ol5yhpy3OIV95Pg74
nwB6oV8CupTjOc9jkoTGF8EVuApKS1/7QmjInaaboQzcLt39TLOsaevO/1Cflw7K5IhA5XkSu/dx
8lMzY6UqAjxhnX4a+heKK1HYjUuWnZg4g6tGgtw3djXl+F7hZYa6psX5WYx9/A8kQZkHpTs5sYhR
hn/AUIaaZ0/88cT5qFEoDqK1d1mNYGMPtLG32cYt6j7eyhQQWEctwQu4StAV0qHdkYWcbu2eKUPb
hBUMgZnu6OWnhT9Y5uhvnBKvmXNfWni51gnugE9u/9AEYp8nNTcy3RmXIBKBNogkF9yE7NjXgbhJ
GbEsJN4RAwi/beW8KlBhIQhXAUOzCKY++UptqaalRIjuwBNZSeQIzKRmDSGIZB2etjRxnJW+r4nQ
dmfghwDzP+MF7M1K5BZ+JJhtKy0bOuId5gyVUWX724ZOepsq+GlS0cZrUbak7ITHXe6uX7oU835J
F6Anb9LrRMw+UNH4CArb+Yv+v4JZhRMg8X/dPIN6NACZ11kLaW3vV8LWkiP5CscMQ2Jhob7PqITS
B1H397qRtJbN9rA/x1UlwDY/z+BYXhUAvBvFG3Eftuinu19RvQUIxKY5t5FC938ZgkiTCXwcKSNx
ebQxKg33Xhk5zMPAVLSxlYdRjxrcvcJY+btyQ/PpZl88r3Vkxg+xcwzwo0vffI0Lxyjelw1GKR9V
E88gWE4TSzcILRJuLXKJb2w/QAPun0CeGIQ7Kft3TWW5dGhygXx1cesNG3kkocFhoQXQdjhr3s8N
mkGRL/Wxun0BWY1vjVy/Fdp3R2Evqq5TpGX6GfmXTAx/lJusevn8oVNf+QPnItYpbJYKvLRBcNTv
fJyfMg5oX6WFk+ZVHQ6+/IqubSaJpRzAATsIiIQM10zjyxrCDeQPACmks6ml8Ez3WqXgMmUodkjx
mQWxpddhc08DNgvZS7MElIsQ9995ClqzmRvh9cmU44c9Mtxxk4BddFtjex7n4Jyo1CaKtd2Hz7kv
0UDU3Gu+LWMDASwfO8VS34FE3SCxR8/Pb69Xy3UPQ71KFVcf1b9tskK08oMBH8fVCYORC61UcZYn
0LERlm76YMVRycKzte3t2tDqNFSJO/cluEP8LYMixE8qhQm85awM0W0jY3L5V2o6Pv9mu2wh8qRr
KiVBx57g+blDmWBI0aVn4Exu8CnrRoKh0BsdoYeP1b1H9TiKszmFJLyvUM5P9jffTGwP2qr7GqhH
6r+dhVZhP21vGmpuZpF9hI2UPQGJ/6CZiMVtDK1f/A7aXaNIwr5m8PRFRrkrxWqFYy8dCAlhl9Kg
Auh4olkdIe1XdRd4at0ElGv5HsLlsVPu0ZwNuI0xxdFZTCxv6JuGW8SukyginvltU6sVX6sD2ZCQ
dtxe7tRYa0adGlW3hM9j/4oWOxeiI/9Tx+tWAmZPJJz4aIZ8tg4Wf9eg/9oQP0mtP3iAw9uC5hiY
qKGyUTr+KbvXpLKehHIqDAJBGvhY9EjO1iyuhXrSe/7e6B2Mm5cuAgY/heNumQAciqdRqvFIEPPv
gjgBKkvR7LozDa7EzDNvMEEd/sX6Y7+M3JlhozUI9uZ4mXucyNAaQnqdGnf5Ge45eXEiUjzuyrOI
o94HvQfGNZouNmzyH5rmq1/FFvRuLpuD1YEhuyfc8IDSpbyWpZKyQ/BOiwY1TEgpZ7eoAMQK5Hm3
pwj3T9kHmOqWcl+PEXMf0naDBrRnVGvyKQKIgBNHkajIpWM8oK8ucvafN8Alm7l0yxUmC0xJHBlt
VWz9e13NdrsJWJKo7x9Q4y3c11WAfxK7cUWbg3FTNsoQ+hO+lNW+6YpO6eI1KJm5hfriEZqBBQ34
jOSsp/HRVOdyfp24c9gs1fSKJzfbv1ceO7icoKppFFDV4QMjsQcQtxx/kPwkofTAf+ftn+p8i/1g
Y8SkcqZpLYxq9ygFWO2g3/jLljPmw5USdPmXczGOriGZe3JCjBlTHLN+NP/7nh2wM/YvYtEGCxXX
Qpc1G7RthI2cWu3NZsmYgH4VUJu3oCMuNv0g9Q6YCH01qtz/HTAfj6zFGJ3LbFATTh5cl61+JddA
gk4sxcK/6S7qd59pv54D9dBy24keYzPfBwqT32ERHr0MG96Q7KPr8Mb+O//te0l2s5HpL4ovkl7q
RrRdke11/maS7pEsjlDhYdbTdsih5l8cQFgz2oSN2AcBeLnM9kK2VaZpwZFLFtsVvIh5n6kFa93w
9mMJOpZGE/E42RcSFRJ53uFCLNebIUy7/JHnWD1vxyJbhSCH6hEu9PWVTl0pcYOPuzUMhkswjO5I
MTNwCF4/XqGKwm6f0f+J4awMOLI8I18rZDlU1biIJWCS3WxAutULObTLe3fKo7LFUtRM34/UOOcn
W8w4dgvw2gmaQiVy26NdSZiScgbw5W0sleIrO7/+bUMI2huhbiuohMk6HZn6oXxfEr6ngCfcrkhW
C6O3qcIN0E4n9TtpxIcmlQBfBHI2wV53pTm4UakoJhfH4yyXI0QBn3UZWNNUWtOh4ZjZ7db2swgB
62t5VvqCqmggpwSdAqHMLVuqgepeo8vmpOlP0MBRHYgam9q4tzLSTrHevFVoSvjad4jsirNEbQXP
7wG6AlQj5WVWlUXxBoVHE3eqEsbv3nOYQ8bwwRKPwMuy+0KvSg2pJ8dHkUcM1lTcvyePHSdYrlor
Qpv7O1eN2rFQN/EKBOAfkI+hZDI7oYmzpjArDxmaeCVirA1RO0yMElC8G/cM+d6u6s8csuzkNxbA
mGkm+YGydRC8GAEISoPzoQozqG9GL736/jLzaodOyVUskgZpdejYEAgivqStIS17FeijyCSEe0z2
Vtls4nT3aX1xKzhdEc9HFW+a2wWEPYdGzMSwhe3DUeF6Na6OOYOJcX4z40apVgfad1yxlkrHY3SP
u8Z+AbKq7kp8Wc5uetEXiQlFKUg1t9d3vrRNRa4+UiHjqUDRVp9BHax5n/9kcrY+KShlyI5MbaZZ
F31q/FCKPOcUvtWRRSjM843yIrW6q4Y5zLwPHYhLS1lXFwj6aq6b6PUwOoBpAIbXuDEyP+LLnzZI
ScMAru0sCN4zV8vPQinLfwgB8kRGcqnur2PnaMUUobcOMNjB4bn4zRkBI+ZOi2eXiLrvlqPZTP4m
h0rK2adQtACD1g9NGb7gpcGKEqT97eHsdunlvOHN6xYLgdT5TT583CYyQuKePLVA+FQm48L83jmq
plfGHs2/9ncYBhy0MTRLTCJ2vSkHtOKFRayGAsSupwcV60tFvYTqxw+szAlbauBFtJ5soDZBMOfU
4tQVIxAfvrCYo0Z3dVl82sqKsKt5xEhka1Ecq8rYujRaJTnfFs1jcX2nAOWHayNlc14hqOJ3Gyld
qbjBvVUd/3TLJo6/wPsyKgdLyDdXMqfq/eBnODgNDpi+X4QWCm+yCjvqG7ZxIK58vnMZBK0WeJDK
Hwi4oGrZItyIzkus+rA4oCBGtGqK5wW3218bTHoiXKb/0G4MavjAieY2FZ8lsDiD7L56E/TPzy+6
QMGRxD4teLMXPchsoXtOXg56mfNp5DYNnzklF43GA13wuyLDtukBQY/crpczOMxd/ROf4rScPDxi
1jRRdiqwOoZRRY0OIxHAGkrGXdUj2Ium5EdtkOZHyS01PpAAfFJkOK2hYAbcTQ+x5CpVDHvByoly
L2NOy4PwvOh1QsM7isnDyke54FZkeNlohbbVICl7KtUkA1TabS20qujBl0ovSRJfSh7GKEgx6JOz
2BRGAHIXWfPdP2rLutJ0qgfTEW3i0+s9pJNNlk6bMlA5nKf5whVXPsePxn/uwIuvqBHj9WdQ9jTJ
/SYA/rp7fWbctCCmCUuL0tnuRmPh7n3FqRFR7dgp45LdD3binZ6ULQvgDs8q9BOyRSlqKU3lGhSf
DJjPkKJ0kZBw6nTOPlp83AP6xquylfXAGtXYHBNmDJjTQg3o2eXarnVWQnZaZNCZ9r7h/AAztl36
XBIIJE9piUb07cAosSJk6z5/Bpsi76xb4pjJs3IbaqXE1Ss+1LXlVOnbUEmYv4AMQoPzf6a+d4tu
lt3hOUCuX5WvNofa6EvFrI06flkPWnkFIJM5pwoiVDNwLH/44l7dqUnZRzeNJTe3uv43Bw/GN7uv
+tpXZW2QjBo7luPwf7NE0WEG+wcfSrVKRQUNo1qP6Vl3I80r8YHWAuRD0DohItEdpVLvM7LSuvYa
RUzmBiwJ2iVF1/bNqboHmxIVV0zmd5hleCBH1dYZl7Vqy5WkiEOXmLnWKE/eU1pGs46XtcC9J6Xp
nEQzdNyUOun0eR6DE5PbN6Q+S0kljihKrN2pC1zDdNkfVaMSYjupHoOt8VuDFH71+js/dK83vxpH
dya64izMYRjMtnYUG/FgxGeHZYFZ22guQe45+8dSNiX2P88u9WXJ6J5c1MEXnjQN3Y2IskO9N3Rn
/fCqrbhS88+R7IptzLXyus5H+LeOspL+4nEHxTusEb5Z12S+jAM61NnEgvRI5YLcNYVl1pdLkvUc
XO7C4GWVuSbhyViZmGcfn5FJ2LcKPO0AnD4wu+gHIRNiz3zvbDX8YiBiThBgRDVeapgm/TaDGMDb
6EZzle8if1HSSUOEuEvhLO7ER1VL1zV2yLVfh69RLyvKdpAX19I3myqbWv/rV+3ye2d9Uu6E9079
hYaGUqPZcvsRKvaQ6wYiMo6xiqfesPa4x7xCrBXMxaBzWeqk0MAesRDOMHk2622ugjFb5CEotpJ7
//6E2/D2cLvG2YepNtwLnXNP6bvbHH13jNmORLzUk/vKUBmo1J6GiIocqwp8zYrNCUtzEZUKBMxj
xXd3oLBbGe0rdDel/5Mkh+62Bd6XozVfrLdKwITqUpQd7t5+rjh3EEEGMV3TiOXdSMdQk7tFdmYI
dHAwdYKd1JO1yMGyNqtW2aVptFbXRuJ/JpPuafooBNGKanGoWE4dp9+ShxxDzdf8ODXWD2gZLS+b
Cbn/ZLAqPWi02/5KOPdIEZ/ADQyFqHx8IYSiE++KQ0rG8asIx2vQJVtpuH+nqKeuEe90FE8hooNV
csGlgUuyhdQXmwi7KiZSga5hTsR/j3R1EZp2jYknufocxgsXy2DB0Rmmcl7mYiC21xz3Rd8XnK/G
5BNVrXpwVzK1mJBKXOnyFn+leJUyKqsvzxCVpzoGf8S5TX/j0cL44H0yDj8Ymkn4D3+5pwAxxvHW
lzCX8q+NCtq4oivzLVpr1jLxEfGZdV/raQSf8BdYEWkW9Jeb69lcwJQ4/x5doU2skSoyvnkliDo2
xrQ6HlLH0YSqyNq+Hf7+alJjX1iqYvU77RSxFfxcwMHegnYJZZpVLFe5xsalnWz5FTvbtZIUh3IA
KZRCREUsrkGHZ9t3+fTUYTLMww2r/1EDnBFiT1ZQtTlfLmi87Bw/rO3EUNhqdRbnkDOENfCBH32C
ksVDLgvIPrMWLhoszIo9TVrpHpM14rodqKz8Sim3N6iDvZCV4cDQds2H9/XRZdnay1R363oMKV7g
p7ACRB7P2/p4d9pip8luNTc2lPD4Q4HU3xTzHVdi/neHaHtQvGOCAtQnY/e+eeqs8/YPHPTAhaBT
cC0MnZXFHJQsxuFhhBUmUDmsbH8Ut26QWaZ9M5qS4uWdsQN5wT0eOtvktYHiZnuxITsMDxTdAbI+
gJz3i0P5MAixbAxaP9SK9hJywYZrTONheOtx8qskYSfCJpsUabIrv7FfEanM+acpL1BxvAtW1SB2
SUyY2TVtDP2PBd/2YQNp1XinYEoTxPE4YcAIzU4cjZ5C8wdnwA4S/lsV05lQ2ZvemYFvhhYR2VJN
vijcilv5rSJ1RgY6z/OaQAngUi9OKAx+70TpkgGY3s0+yn38b6XD97dMV39mGxQWUCjmy3Xmp8bS
T2ksjqLmvCyvJDLOz4BacVG5N+s+xkIhJACKTcgI6Gvd3pqRzp9sH4OynhKLMF2REReu0hz7PmVw
GVUg0VV4G0hwbAh/WUH1+8R4UWDD2W2dYo/zVWtFUE3fa32GpLwN1QX4zoQAuuLva+ynLTw7A337
TtY8bPgFlLaHzH1hw1oo+nBsK5DYFOzNH9774YfnaYTXnvmJUKkUpMONSKxuJ3vSHM5BgUwpKKgg
qkbi3dxyigsiEPw/X8eOPaUZwwkjgjmDvqRyzx/Z6WUtbFb/k1W3WEOYU4T62inlYSCqaE1W1DPQ
NTSxbsuV673s6rbTUkCjXu0sYwwIDhEX+atDGTU3lsHb42mO+24nYW9fMDvDpC6JRPfiZFzflcLN
9AzaGxefSEnww8HWbIO1F791XUcPbyUWU9vZ9mUJzSysgsOauGGXGLOeBXeRqcALhT5E61uQSmSt
7nZ6iV6Sbaep3ORZHIg+y7nw1IGkfJeSnCzrt9eNthpbZsSOlRil5wy0xG68AN9rx6nm36wg/fwy
s+gJfOHyeRHJH+ZqZLCXIcXCAmIPJpBkaVmauDDcqIn6rQkDpS7AELGz1Ic6HC7rRhZp2oCcGtv5
zjzEsw3VloOWXKWNzWwLNFJRDYKD9OQeJU/9qNqqCyfIz4RsWdqNozx1POuZb2Bu7X/vIfPD4S2m
WUyEBEFA7rwTGpmYBsrFMTbfXvmN+CRYnAybHInDky8pCLD5NCFltNSGdHj687k7Zez/j0kuWpgR
XLBl10aN1vauKIjy09FXvAekR564ZKwOY/A575tnVqiR6ouUI99xZlM9K5WVaOZ2PwKggLxFsjoj
g4Nte5KR2EEHcM7xsG70fjJEEyu0qDrYB8K8cXGg1TQFzrGYRJIq7J9gzVBzwUBxjgo43AXFD5V5
DAWlZ7elWV46hCJw/WxTs5QtN8PINmAUu103VGkWTCXvle1/+KZbgTaOlhT+i1hUMFF/hk+1BBH4
PEUm/PHbVTnvPJ+FK1r5POJLrYKWBnhgMkCI4nFeys7QD28gkbnH5Ezsz196MG9HC214eJTSJRWi
hYaswl8napO1k2e/hMNAn0F6hgg6sU1b/4YAReh2SmeUNMHpvOs4zEnwEV4EzrnbH7Bky06xQ0Mn
bk7qTOsfvVkIgn+I3mAzF3kSoM541//fmGuqDbqX4mKWQ5cQxaJleZ722XWVkZXW2Ub4Em/IkO3+
+PVdcSBuj4SkopBMOwkjZqgC3oBUO28JEiYAoz3AeVeYOv8Z2lPkETYQ4CRQmfSdoYbzAKodUVuz
IqKmk5NZaDXf2Z8SO+Y0bg8TerL9L63HxIfWyegLIhjuTpkrEnRYEbKNU5ha0b3bNGipLXfNes0L
7DhSjK4nK81Ky9ep2xGqBNg8EyaX8Tlo6aQaAfZX2b6bRAfZJ5ZJyG5geKr0LG9xNSEotOYrgQHI
N15bq/PcbqPos/uPmkQUqdbc6U2FHmUlLCb9EER8C7gA8Ddpni9r9FlUoZLlTPkSRyNnGkipqfhV
+9lvun4DiWtpTmwvykQkKdVz4Yf4G40NHcrMVa+Rzm6FbSihS2os5uDBY1ceJsGgoinCINnvvngB
tBo1laHU2w6CQd+h0eXH7tPFuk7GubQREsu3UstpRZxwDWkSojhPlQltS6LVzCIC+Egj3Gv2CHpD
Hsvf49LZ8AbiW2+6EYLo2eHPRLQV23UPgliJ09E9eLcLOvIV5xLcHzmxXJ1pBgaBGn7+Srdbx8WR
nEfjr27tuRQxFKj2ijM/ADdXXjwBvTZj2ozCR3I0mQAW264FXaHUfY6h+c1NtcRbc+Ue+mAijOXh
At1BgXDN9eoYk6HgNjJRMAaKe7QzfuzeLaK2fRH1cTt5ALMM1TBBwqxO8bEszX/q1zppmh+f/Qpv
1J3lGturhU0Sz0I5ClTso23ycpW9WehYuaxqdwwq0iyM173zuC1gRCoDGYDIh/QIczGX8Er3mGe5
OQtMMH1uaTB5lzz+CUy/4vxGuAHEUOJzSsNRhOfGtuhy8CzkCMhtlSc/9ZD23t1jRD9BeASdMFxK
sJICQEqaHzh8e71zorAIfaUrXFq6BQxUSi0eg+bnMMRp0oJ7SsAGe1NDhqVomQiJt0r1Rg+VJNQZ
PyuQucdLZwfHZmlzf7xI2PxGdY3B5mEoqK1byD3vmJS/CE2gq7NhYRkQk79YXuQLqxMIhSEiwPp5
9qn4K91PXuXnsXwAaHdG+d0H5PYUgcKtJJGl0c/Wxs9l5KPqBNKoHbu/7dQMqLmLyw5VS8WtdG6y
feB+Tso5DeTEIIWjPBBorm7D9oz+WVVXxsnmnbymKIX61O2qYgF8DrQCaYDiab7SERJjwjmEBgJT
UE96QVD1RkiPuRQKfpjt9Z15JbnKbV9hSG9Z6mCVuHJEFjiNFg1CCcCEuTxPXh6tsF41Q2pYqtT2
6NtinuG25YDczhZv2lTKzg800NkQ5m2F1l4peDiLuSBQfCOjka362yIjlJ7Vt1M5W65qGowGdGlz
fZU7OPWbnVThbWUBheTIWB8wJ0SPC7AjUAC49tQtas+kkjrN07Ve9/WDBetnUwCQIkinEDAlz+j3
8WSANekn/J00TLmW0QK16wlKs7LVWAbyggxBrVGMozd2XWYnzeDeuEDfsSkAy43dG0ifgnHuq9W1
vz6ULDtUmcgGXGTD7kAcV66otmjSt/mvcuh9iLm/JVT+XM3KtP/KnYUchRu9Pe/75dik/NAfma3g
eVvqn1+Hu3G6XLUEr5yTdzzFG6YrlipnFr9eNYHxgnF2nmpTKxND2Pf4PiPrS28b4vR3nro5yvhn
iW8enH6hqfBsDMgety3Hnh4v4qbf9ldGi6LIHDZ0Wzq28WyBpAIE0RmMOhUdxSOtOWu8sfUC4Dp8
jMFuekx4q8OqNMCCIO3edTqcc4GvjT1MEr1iSZMqwLiSK23XOy0ryQjxamOhj8IDbqT1vEN/LEvR
PKasByQxq2+5gNElvqPP4iMZUsz/nkZFdEVFb+lc94BKb8rX07mNe+EHP0n1vv7f+AhNAB0IC0n3
9IhjZIi4CBlZQuym/aPRnO2HoL30V7Lo5FikAmLRe1pQZ2q/V72hUH1Ce0fNp5TB3FfbE/2J4cxo
sW6jdxMTTk7zjBKu6M7Gb87+R6RAInSB56p78FsvjMDqknu0YJ8e5Yt9CQAPQf37thEK7lI4Q117
Q0q7F4V/fIHFn3yRNa8HYGlxcRDVoa46F5vnETojnYbrqPIvNit3gwYYNppzM0+lQVH9/GDpy0Oc
ACZ5TDAI0uBbPuNVQ5zLrH8bhSiQURbwQ4Qu0ep08rA4UawsHcV9LO7iBEnU523WPGex7+0c1ICT
Q0LCd0yOJKuNJhElSmwPKOVu8Kv4iUlcyduUPwcIfXdMl5ay1oMLkSSRm1OscysFwjkeaSOr4kMm
iI0MVSdXLzgAtsN0YIOSdbhxHT5l8MdqIrdYTMm5pZsIbEZn2303rqWWqQ0JKIPN/0Ox/jepmRvC
un7KgMo5uqpSv9Nw0jwfkhczLonUMHkefBqjXKRpTdc9ytkZEWzEHVGWl0t1SsB3Lb4mmeJ06PES
0l1Ml2e+GdO03xDYCLVdCkOmiQD0e5kVwJVa8LhsmiD/iJ9e2OpYglpvB+AmQUzIT5RWgykJX7R1
tPZm6x7fv1zBFB6MCP9mSQ+yUat4832BeoB2+QFY3yMX05bcZEN6bp5cCSyTRvYqOybJ4mw/gbLh
k0QjeHIO5+GAgjvpYOFF82WUoSa8eYdIL/ZojEQHOlqne3DV8L4VbkNHWkCLm8aTy9mxQUYdQ20R
/Ld6V7HXj5r0zd5ewBexS2CXnIDJqA+Y1uaNdcpEed8hmHX3UTMFUq+eFhaGFUXUv2P1qGRDtwna
HzSKIv+hfoYp/mnYnDAQZScy+7KfxMxaxP+p5AGdSp0ZWsELDtsuiYg9/beg+WfHuRYsxTqEOEgO
dyddokpE6BPu9EjUBNRMCv0cSdR+28t2B3WFr27ooJJGCkK+DWfFUSj3qFpge5KKVmZ0AsTKzawW
j5lMEjmssbmuVmENgXVRLAeBAH4XmZYOIvzCnxqQc4Unl/TmthpRp/v3EiYc1CFmUwmb3C3XbHrl
O47IuaABX8DKg9zVFO/ztcT2Nvl9PZnSLuWDt/3UO7zVT8yjIrhVLcfuta5u6NWH1EOFQPkbXF3y
NaGQZ6oGzlUvJcTE7RX6poYqmlQ/EyOyPZMMkpcREFn5T2biBE6jOVHwO3B7vuugEQSESuWgLcFS
eUaz0YP/HTocs5yJBkkPq6LS1fTOmMa9H1vUVyXY84N114r/GnArO4FBAtbsfXXhdYLlkRSLyniX
dmqf06GaxeRC7vzvBbvRYDtyoVaSJNCZVm2aegEUmhbrZalPWt5mwj8CxsyikXwrlodJ6S9vekKa
w0CxB91LSJQbknXdJzJ/o1Dd+jWphLKWOLNimbxeFu8t6yu04szKwfMQjd+eMnh1BZ1eIc74FNrz
WYBzTD+esKjjc4CLh3JfyFqsSTvC4kGiMa4iFU8WpuKp7q6r/i/IRA/4fxA2z1Wrcng9uA+N1ek+
o6LlMk88TRe4srioOBXTCyHZQgEVRf+QVcF+lJYXCTcjz4XS9kUAqOolhuskcBw1zY0RXqviEGI/
AYhOjE6CqzHvlRKo/B9/vV0dml930VcxzRPSeY/NEEtJrFC1NKVfg8JV0gYE6UZf/oQgkBQJO0lQ
8J/PxaFpqar5L+HRZuQ1QjYD6CwzQ4+1QrvsAiyPKz9QVXvPV+CVX8X4d/xu9fG5BwyHIk4cYTUp
P4p5DinyiykqQIlc+UeOPMV2Rhf1RWwGS9Hcq5O+N2rJnUK1KFxMJJdD2I9FRjW9vtWc0nZLr6Ph
iKWsq1yvd/5Ltj64uQm4F/ET8dRN9cTWFdvw/6FVOc8mQLEK+4RTRaUPKFfYoqBQIqDF+s0qUpce
/5/XJpUT1iM3viVtUGqKk/myJT91FC98RMPL6rmBKhU8IsGN1Y7KfLPkWz5IbDcAvHNYyjefFqE0
o25Pj2EBbwou1riiuD7GWXwBfAeZ71d2l4TCA+tWCWD9gvIG5U19nvPCCmf5v4rTIXLP3YA86sO1
8+YQMqMdps5LQRxMA7+5UC3OX6f1gfOdRJEXBl+OfpvPFsHgowicpnIsQ1tkezL6kilaCM0a1X5k
VGsB4NqL47V6+CMLrV1fLqcBJAV0lEVmidzzIbpL5enqOebqRaqU01JXMcSuHMlz4hc3hN/lT2+O
b/ZyqjQDkAxRCg7D07PgPXWYOCrVJWXE/E1DvkuKrvmNajITxrIcyCPyOUEkpzoqpTJEcyY4ZIBd
grZMbiLUUNY1+CL6FfLqQ24Jqvog0wkUdrr3sluCB7kGbBp95GpJ/Fw8w8jWbK4S7DuDHhyn7+Wy
1D4zVG53My3a/QRy1a5EIDpTy7AO2g+UatXpo9P+GZIZfElWljDcJfSO00qf+URB59X8oA05z1eB
cV40+uW+ZK9taLVmKlORk8sNZvogIvz2pupFBEMef9NwBDlWKRM1Dg8CwHLW7UKMEKesuwRx/uic
hPJeHq1frR631fi1vXXL+3+0dkz11m+Ppr5Ty47LucG9qqRZ4lpk5ArKCEcBNC0802ct7y5KsGQG
kXyukK4arx525s6uoojEWEZU7PSN0uVwVQfEk9WZbiOTwnXljHrDoDtVRBpgNVQ/+SZR2MBvevqH
E7M96e7jiinEfXMLs7XHlpEVo0ER0FunhleJ+rZCdxheeweWLQyoSDz+w/v9fkBa+V/G0QgzBhTv
UDD8RpTQtglw6UCQN7aFyegQI+7oC69TN4JFwAeuf4Yl0VdADGIl1vSGvcc5rWYdLl6EEwrECo2a
76QW8b2umU1201bBP360CDMEzsxcJhUGIgQ//yOHjHG8U7bUihJTTe7SF0JnhqyBg58ShY7PDxOy
kz7pz0oS6fNG+HqcOy+Hl8f9GSc5KauGzwM6A3cj7UHyC73ao2U9/65Or/qjjhTm65IwiVmPQazP
9IziDZXVmSUIZQS4eQ0i5+CllLQGPCCRlraMdzNU7Lb1ZD8iQVsFMnT3TrqxJd2PshU5TTryxbaf
rVYKfyYEaZ9PaDrFOC5zJoKb4xc1zNffAuMUGCC//tMhm/acPe+qA3yVPSbs3B1db4DoN41Z5dG9
erhet0lits2z/hc2MAnUqmLFxrMr85eCpcp2YvswswAU19XfwTHH+TR61H12BAUOadXVDy9hf7z8
TnQhWjY2eR3K2CL3PRsuLeHoPnGZBYYgNZTMYuaoYw1XbCMqTTYSX1UVFkgI+fa/SGp3WsrHxj2z
5GNoIhRuSZQFl/0AM0Itgead9ZhPmctbcFLmYYQiiO6mOC+jVbiLXumZclZtdMuM0E7z2kJGoG0T
xBtlMATtE0c+uljXyIxplv9vTQ59ncSaj1NUMzb7wVyXe5hgBPPFfFKnvr28SyqnLC2K6miE+L2B
2wQ/4FypSVMtlp5IxFVNfar9SmXsgVDcOsLsWwezv4xHkYqhZ+PRRVOGbbzBAjcclo7vZhzNfkI1
ynqqH+c06RC5nnAOXxzRchoyAqFnAgbpXrgf1YnFZGrVfg5cl88SJi+fO73ieSasHO+0fRnLkOOd
J5VVAscPoqkT/heziG/D+UE/LpOob4q2gm+i5tjFTGU0rwa1HRjTHKTQ4dZzK+ny2BBkujTIIGFg
UFJw74EEVsnAtMMQ8gIeHzyPUAgXYu6R/CxsWsAxZYkbXezCNe7Quv2P4SOvc005Pvv4f0Ci/BZZ
ccA1DVw9d4I2Tlxm9wVDUwyk9JHyqQsjDKG//KyvkdK0jJvZUHhNE2wmtNpQTxPHw3ggT7AqtgIm
IZ5VufzuWXACxau15bbiURZi57S6a8jse8fv3yUfCcmDKNAsjvY6EhjVWB4wR+3nB1/6K0eMkyHG
MsIJOsoXVF4veK7nptfzO5mgoVgphOUO+Os1/Pj4BYC0nkK2B8YNDfdNMFwCyuHh4pZOw9FpZ9kW
2A+ZbKbgujWVpIA0ZL8PS3QhYDPwxiiNfGQC4rFA1ReO6pRrWt6x/w4ob6YRrFlxMEsIyYPDM4rG
vX+hecREvJJMtup4OTpqOdTp5N35GBCY8akDGcKM4F+grXFfKTDrNt1tZmggM1DicOozKjBYZQCo
eGA5QZXc3Kc/NCoh4d99Zu7Utja0bPobdMQSU+wiNhn8f7NCugYgYIUaJqacbbHt23DO0puEpDgV
qth26B4pGp78ZJKXVF8vpDhS6Fga1t4y4JKI+EyVPO/ygLtyCbK6YY3ujEThUriiVQd6Ky11mpYV
zGyDvgGY3hU4nHuMBuWvqCE1SJfgXloGKlFaeiTqRmLbqgTb8+CqrUKxmi2OyE1LfiPQrMithS1H
wO2PzsxHcDp7oRdeQnr+vSzapUc3qpv6mPonDkMFjExhcV3Qd191D0s/Xa82naYh47y3gYDthPLU
pFJB7r1yp3xBoamtJZwiwr/3ru0LxGgqNld9PDPSW5JQFG6jcz8I1lf+dhNYW+h8wQ9EtkOttfMc
Pw5iXiCcTYyyCGIklcZp1F8Xk0+LNtikF10rq2GyO5YMQ7t0uaNARDHgbBPS5FaQi+cPkO130HtT
7NvEVtnZ4ls9P7wie3xnvf1buLHV8DlF20WX6gOBCrtSB5S+Nfwtf5WR8kzyURE0c594a9SKrVRk
4JcCC+8wbzu5Eqd426ZdVZIP7w/RL40dhCAtym8M4yhItIBETZ5SlxdaVXOfWj/lxyDl6Qnhh6se
lZZkVXoBTRRW6/4SpiyZLBRC2Vi1YO483YFJI6UmmcD3zyAmGWJHenW28pQFyII8e6LiS3r2nAj+
uSQ/Wi9PnF4ajB0Jnnf8MhlnZy2dk7JMcddCRhl1GyXGJHU4PKOlwplLXhe8D0XqiqIHYV4w09w5
RFa7E1WAMIaxM+APG9vv3wRiolz9+4HHEfUekBVUOdkHNg536UN1oh/CL2pjRUqdHRji2pRacB5q
bOKPVT093v86tQxy+zDei3HP5ykUa+ZhvrmV++MQLr5eFlqx0IKmwQMYspsC809BLEglnytLlha2
gxuD/88fI2jI0gMQ0Uaen4zTRIAtbv5Tqo70zngSkB/JHQU69h3Vr/io/rfwCAOLtVk6YDjwxVdE
f+lGPkYjY4Xy2ymEDdG7fmJrHTwUxgkderRTOwGF9RRbIiMbOR7UxgLPl/D39xeLKoWIg/iLvOzP
GrZ7CPmrfRtj3O2iL01SJWMyZ3N5icmU9Ovo6gqK1LQalPjbnAZuiHPTEcFgCozWHZQk/PSqzS+X
foberZ+h8gb5iRH8I6yo598nN68+Qhe8mOKS4LmvFT5ktNSvceTlEEBHILzSqwmWI6PjnvRdb1RH
Uj35KI62rYkry919HdZ8BrQgdgoSOPzlBP9y2QcSVTgRFXMOSznPzNRlQEUrPrxo3ZeFq0zV7YeQ
/rr0IgjITK1Y6c9yP2VhhG4OtiXd6ACdx2utYWkB3NgMGFGVHW6GygEq3PLG2oJ75qHB+XBhB+Zy
Sr7SMxIH2+ygOeR0dxUI6P9gShNGyek7cseL0B1C7sZpuzu9ZTjv28kGxL0OPvP//xeP46ufrpOh
Grf3M14/7qGUKKJcQkhawPwi/i+Upf6mk59ZypX5pErgqrGqhVLYPe6gK4/SYRO+HJzKURr/orNe
fsOUBPbQVjVM7ajqCWIkkj7tRfY5lQ6DneVQL10u9WhGXteLuXaB87yRKCxbXAh4oH/LmKPOn+6B
LRktLSJOfmWEAUJctkBeqsZmBQ7Xkt7ZOwNQrN3ZedP/BZIe58/QDBpOF1O4uVHFttGH3o3mJjUG
Wap9VkCum+ZIy95fP0gfaqhYwnhgdvn4PSh1tTc2KpQbbRweB4a+chas7BCU5vAHjqsDC99zhb8w
xXBUVGzCT6SfI2tnbAd4SRd8jiCD+SKUn8AKgLmJHWmeT1RVT9EuMiijFMHjpzMQNIGN80LHA0SX
hfpFNEPjcnr3dNMsUcA68lSi3SjozrUTPODN4i46WHjuqO0GyBHR9AEf+QX3Pw45bjLictOoFI5V
ZHXwAr+pqLYqQvwKig4b4iBQbWOvb4Ukj/jp82Rn1Mj2M1xtb2pNS/OdLT2tBgw7HHZeGS3JfwOL
3we3AqCQgHNY+hMLrkxQ/43USloSomCNPxbg5ImynGh0qXcBepSGuorcD+0fNZxPwGL0hqOfkpXN
QcRVRZ3M74f9YZHs4py7tquWXkBMYfgrHwyJv1rVGkEKE6GHCOLAjUkBowjYM/llZxF6k2Roli7X
Pwqwt8c4m4M4ABR6+IkQxi64/+WGF4QAbFLxiV5I7PbyLT8SDkyAKAfX/GnQJTIVJO5Q1kFkbmvQ
+4p+CJEsgAQkn2GxYOU4LjiUWI1w09XL992s7XJFdMn/jcFyNPSNpWGS2v60SmVm8pRm0lqpU22W
sQ0qjTMN5l7UdTedYLclt9JGiS3cBRFZG5vUfXfzsyMgYuW3DM6RNezemiaBxeh4E7sOcTR1L7y6
RKCKU1iQLs+OlQZNnsHxOMOWc8Gad1DhuX506eQ4cUFde0l3m0t1ZerTVlf5tw3tXRyR3lUA2PEm
9M6EnJmRZEhxaJmw+PkxtnZiDZITABYD2zzWlDseuP/nOIaXdbE4R6ZrjCLQjct4FnFhgSnB8mLB
zn3KFW3DiOHuEuWAXEQ7mhrt5WSducUvJdGxnkE9o2AEG8PAnhAPKe4pEKfSPKJamk4ciBjwCiNO
403TN1tNxzHiA2JBFZoTKhYZtqiwXT+Rd07YEDZ2ZiJKWfrOX1TDreQXpESFClODKeIOXHNReat2
hz4qLusJB6kh0eRKX/czKRunwCUY17cqVw+cT+6VSEAqoxiJ2ubJnrZk2xmWWlP0EVFYzX6I7E+8
XaMs+IBShSNXOrWn/njEGOu+84E+GVPWgnylpD/1x3v3KjYL+iMuiNSpn5w+4/xbxGAkStTF1a8g
Nzp2HocgIsUPEjDCgVDLtwTephVtvFX0s0+lBSSXG2r2mFsWrWgEG+WPW0fbZ93A6p/4TX2UHf22
4Em/g8DftnjyhvSXQPj3ppinRLRzsw3Olirmn8kapyX7zuo7ARGhumdq1qRezHleebcwlndCP6sH
1XhZjoJ5O0l1kCvWLMaNFqVUxK1TO6Rn3QdKnzI5q48PRSgCd7OVlGTEN7E+ACjW3wSJDWh3ZzaJ
XsNbgT+BfbY4K+NBn5+XyaEX9+FVAYlK+U5f4njeB28orVajJEHbTjnig+vbCWobQgK5awVTTWS+
+mxuA/Prj3/8u2RJL0Didj2zntqkkXpSuTvj+LfOXTlKw/DiqPZYfxI2d9b/WVbZdccZ8sy7Wz4T
Muz+WmSufC9kT3ZvPlNZKcpZaDM8RrBb/eRSxw169T9c/NksPgreLW+ylLmLdp/vCI1nNrgafBsh
MRC5OzHy877m/bIMZlWQQll4dcrtdroUaAuM50CYwTOHWzUmtAfkX2VbGfFOTiNT8g/mI45WZNXN
u5qf7bT+Ng2qrwMQUxR9Qu8lxmWQ8sDi8A5l2xE7V4IVvoxP2DgkeQZ+ltkjvPIigA7iJvYis0os
iyn1Z4eRyEep9LCO/944eStf8mM2X0nZzA2Ghqcyr23+s8jd41nvR663JDsa2AMev2wJffz2VfoL
xmo/1aGi2Jwg8DeEfBZ5PLlb+qwDQxfggdytg/do4Y/GEuPdtIu50moMR88p80unRP6Lqlv3s6Lg
5wgq3SPxFDm0p06AY+Gv3tvfzLqvFS35FH1dlh8LAwklrA/ajssoy/Vae5AAyO7RwBjg1a3ew0Zz
V+10DwNt9xeSW0fOYpvkNzyPu5QAWSYNNkiYJNk4/lI7rqXB68jKhu2vaA9FL81Ouls2Rmd2Swkh
LlWTF4CQXwWygbIZKPd7vPm4Hq5Zqr56rcoiyHbmqT62J2cohqZNfl9Kbxfck6rCiM0iZcMk5b7f
TAjUiSawUO8taQi1aAHSwr2ddYQd4kMqFJfUd2j+BhgBI+FYuIJXuNHIMbrIOAba2ngpHyBHdC8q
l3i3G8IBTfH41sVwNq1nd2m0QmgIW/AGJe7jIKaCxXyXlSsvZly5lj+z1/CKUX7oOZmu8o/fL0ge
lJoa4GZsRFQD3UHZsSchPNVrKOELA0c/duemRqhJxGC4uDBNeyh2FNZhUOmPjfs4VXpEI2dmfGr6
tb5nfo8G/C+uAeiDz1VdCmPX4gqTA+X5nimqlWeQzzJMWd66IR9Y/ap3uzJJZFzSq2BcViUJBxPC
tYFcRW5fBEMrLvrGne82Na1+WTY6tYKZ7kVNwq5ZWEKdRbJqS2HPyHUgAO1IBqD/dQOzj8s+yp9V
4/Rg2GWXyzkCJ2ibRMYH+jQJvIz16JaGl6mjOr1Ai33SbMrtz/9vVw0VsC3O+on+0cxe/hoKm1/3
aA15P4GbSc7JHMLwaPQNqjvApHG3Yv9y1OtrMUKnx1uLSZZPdUc4FZ2aMHan1wiFnmn6cmyiEAQD
e5xXUkZcC/rpFDoxEM83Va5HMXVqQsriQm30PW51hPVEQTu/+XoOvXsltvGi3q1WkgWDyViT+qJ9
cE5QKeNMAzlpya39L/lcLS04TT7T3+aLp/DxhdETC1dIuCpBd8S80i9IocqjYWSNv/2fsfyN0XgT
wkGWyYbwuKi2qFq7N4H/cwfYohFttwOpX9aelQavaUj5HujgA2cKxp1Go0+l/2eFOvtZU4yJ9mUU
Z6mmgoVwswwuGuqonb8foXBO9l2rK1T3DvtNfg486koWUlK+W3ZWLOXRg9C4VvlCH38G1MQra7HE
I9CCFIScpOZwD5fJdJJjXmlUZqibH0a7POrESHLfU670eiYWAVgMjjoVoqgW22n0RWHge7MHtnpJ
o20Xi8kKZ+4EdM9BS71k0T5NsRENc3CnQC/os4UW36ZgZBqX2KCpdf/XcO3bMhm79RmjcVwb85vU
eU0zfCEdFuwiyBaNCILclFM1RT8jXjFaMUlXHBS4LX2N6GM0kMS2z0wFbiX4brUBrPH+9DX3g8uf
YzNf26GAT8+ziwmA0h3oKPEM9NgLD8BuoKfAEbjvUzu0k9mif5pgW+jTGPUsc+AhboOq9kbhLxpb
PVIm5S4nuH7OxJTkTVPstfhz23t2nS1RlM0wSBJ+HCgcCADFk+2SbGk1xz4PgLqlBDJKrljU6LE2
Jv3B6JdAv1vcnMYIeb/UUh/SXtqKKe/hTjNMU82bb5/zGIwrdTEymapsOzqyqYCoRYjaXl70StmI
TtH8koKeio5cHmC3lPdC7kCJr5YG5pL33WeIkFktmwtkNiXvMMmQ/IGIOIdTjs+6fsUW/M/HOvRa
pgYr1kFMfdXX6nYtQ9hZT2Pm3XO/0VKMLE/S/c3eCKz00puv6EP6xy1W0iD2MF+Dz6F7UYyH2EgV
JF6doLstkEzegkoiaOZlhq9O8faOFeceNAFic7AK8GrmmD+iFQpgP74BKkdWEfvOl9ogJ3MPCIcQ
NnPvlEVM7CPi2gHOGNHwgF1EN+DFzm3YEAqy+Hr8/+d1PhYEUiofTRMkv1iT6C48t0tT2Pn6KgIE
THJ388agAsig6WM1S+VqATuX2hbnP3G9/oDv5aKDcEaWFHkwLKNSDyYN9U3Fp1+GfoC8dGf9X70C
6ifBoLThf4sTiZQivIzEe4+d4nWdYO+JqB5KMWMnlyc7mR2MmsobC1lHV/FCajdlgPJCUKT7ZIVV
7by1048ELHbcIBODRWIF44N85yKQ0o1K+/NDbcSlT1Q45P6HyPZzr/BUCy+EuXHnJ138dfkjr4w8
GeYUnI7MxGsktG7EFmVRdTjj4XWjhnSJkxJ2WCrYlRE8sgfjcbOyIVXK5NIgPwEC7v5zRsyL+Hf4
goRCjpdDe55tp8qfR5fHAWoi79tp0KvkkTjFh4HKc/fxRW5RubKFSi7B3SggQ97kWDopPLEyd6r9
8R/TTyYc/o0M1bMuvGwatLb9Rgxb+jNAR0w9knFr+Ij5ViTyJGgSccwdKVl/8/4el0aQfO6nkM0B
2Xhjmgw8Spqra59TIVsE3qrbk+yGPb4lm2vqLdbp7wLYYIQVQHV1ZjlGRFPe9jENbsmM+BPbKDLG
1mu96TWNB92nkIWGZn3UzNLOh4OHQI+kR6hfeTrXWwLUkrJu7lutOjnFwDLkoi2C0Fi8Hjxygz9D
NW9aWQJF7a4dY2EkhW9unn4aYaSpjID+GwHBHs4fFuWwIDfLnvbPUnKFmaff9JpJgyS4kZWsX+Ip
LguxRs/75YiPs9Joy/Nsr/RZxBJj/9+kwAwaaHL8zYmjWZinpogoDnjkM681Y7p+k1ZotjPQ/8wy
ACZIa1bt0IlmdwVfW1uRKvwc/PjdprWZ5Uo0z80frLvEQjE48dJ7ukXccY25KdH2PkEZOb/Z1zNL
SXi8GoHng9IXl0+/LTm1o8eCZxhSTGrLfqrLo3yO91B4MrzMhywwEbJdNSLHrJx1X8heNyaJo8Wx
jkEv4UgaN9WGB/jgjGKe+u7BQEvfRQ6WuYidkq5WvjTokwoAq5+lLFV1FqMLMF3FElOfG7ULyIEF
EFbXN4A3dvBcenamPen4wRQE4OUou2hmekGRgBjQvwuXR568g54vXYZFThDc+kaAgJkmnJKPF5YZ
yUsdEiWpeIgdagjnAQ9qL7SWvZ08JC6J7VNDMH7UFaVJ/eJbHM4CZKcAudkHDONyVIFPS1ebbV0a
Ctn11rsMThft49F8Theg76Q/uNHmLsJJ5uM8tuqfBuBLAGJZS5G5mfcoMyiNPF6i4g1/N13qzP9X
hLAY4cDxrRy6xgi0NoZFr0+nxApX4R66Zyk3GVfiX2y9za172X+eahOQOGHLqLszKoJ4WIdq5RRU
xVgGgDnxObTFoLmTm2KDB7Y51iHI8W3vPx0qxK+XKnGlQ2wj9dDPgtinCyKFck9mCIImnNrfYZzd
ueD2yQKhJJX8+VRREZGRAjEzwQ9bZukvkFQ+M7Ynea0qlazjCuhGHTNAuenOuY1eN6icqaxTcrUf
GkBbnfv5/qQv9ufaSkK42KnYXw1Cr2UT52yO/+tWwH6LRyPQW4X8InMhB4Tsw191JfapQUJv6pHT
ksOA396tfbLUf67JzrG9BP/LUJqTdYfOvTmpsxYcXi8Ioa3PmS8FkJKnl0bZpErN1Qo+I0Ob9YBO
QsJ26lecK9jIfoUBFbxPQjDwKDKTWwH07vaq44XyV4GnA9rD/C8AM5cl9Ai5lrBN0gjvDj3qhile
B/mvzBCX9laUTeZSV+nIKkRFOy0R6gronmDaEP3LfmXF7cLHcB5U+KeaDzxzGtIApUKzNYR/Cw2L
hx36RW2wGB28OUMUOWQqTwHx6xRV39VvJ4kGKyeeGME1KuOmd0T0Z/D561clVRG8e+OP2uUjD5io
iQv681FKrNI9BQDEVVixl6+Ddi0TRIbwoS9/TZQ/W+bMklI3hAr9cTUQFfUzQ5dKKJpRo0iNC+8u
QQMCD3EZoohtw6n9oRZDM4aD7IhNxcNGHB5IWsfeuP75dosJSXPu1uKWr7FIBijv3B9yo+CaCmmn
GKq/od5pcdfNbscMAblCcN27RP+ptzREd8vGNFOV8CAgjQLvVcEO+8sJ99SNiIPEaYFDKGAholG7
Y/aWLlGTWzRMy/ndPGs+Vq++3ZxHBruJG0lzOBMTpPviTxl1anakqlHKt+U+jvFNk3H7WsNXpDl/
cIv9NV30EfjiyCcSRVyEaWJKS1blUCS/C8HWWpvBtW5iCSuVils+0R9T0jOHb9cIElaopOzw5NdA
wuZF6WneANXWIDMazrPsvGAaOyTcAwQlE9IQVW1ascv8fDVeH4fnGIhnYVAmFNHeEMCSzRtKSXAo
ZH1JNOlA79Ox+yZPXSXPaTYCVLd2a8aVxG2ZITZTBrLIFqYDzrdvl019EU1iCiZFOhbS+co6nvEW
sJhiyuSwv0nk1uEsd4p1/3eI4d6kAkWqwaYynQlJAG2SMYP0f2D2Atcl0Db+spDuCwF/iyVh5s9b
APxK9sdwZ9g2IoANU3qoKkRKESdL68Dn+vI0eXvQ8aIdrDvkwOl9u8+T0Frr45Mm7BezQzV/H2IL
G/gzkVyziDdysn73ZROxABx1L2MTBW972G2gK0Ur2Vz+vINRTFxJfJwS32kYaFx9gI9odzuRKRvu
lg+akcoqFiw4+/QKYRFKmxWodQ418vBYMBldsD9fhuBMuBm8g5FdrON6tTfMuJ9Ud+73/FVc/DuV
K+oBGn6KDw7Yy4gph1Q75sKm68kGalTI11YLvnb7DdpYt9XwNPD1TyE72Hu83x8dmXYLYEgF+qus
b4+5nHGNChXRgbpP8MrOB8cOWvvutveBfOLsV6vsuJ646EvSEwxnQVn2Qbymge0AlDsflJ5Xiask
ReBocR1jFkDvv3W8NPYJkH6N7ll0yze1mHbcHR9McY8j4mPZEI8PBWXbBOwRUgc73bJ6KqbL6NPw
+Xs8D7CtgJWcFVvIrPyDXOEvgFHqEvZr55v0ilUIcSpHvNK9jfuUz5FZBg96UHjvWq/Qhye6YrBR
QNZFa3+w+nOe/v00km/UnXMAsozG85zbN18A8WneSnDX1ujZkBdSpZZyS3/Pb6NdvcouQN9VqqHJ
t1F/UOuxVEmGbUN+/LjOZDP/T5t1hbey7eZcWNVwaKhIYS+5hdiu3v2c/E76R9jOrI2i8FeHx4NH
Hji7yfleIoYu66Es7fEn/EIjQ1injRcFmR/yBKrIgUVFFILcIk0+cYfDwwYJZLj+BSvRkt3rEIRX
pggicQFvrOanV/5pKi0SILV/BpzZN7U4GWPo3JQoXBfPU2ULj023xNjy9iEZtPbhnQwCMXx11Gkh
rrdBu5Pffqp2kSu91jqgKkr0TWiLyYzgMMFlkU8v4W2wz217+hkTc+hn/9zgv/zfOtDOlj4EyvDG
+FlGMenjdmak3vPzjUAbxndjerzYKcJcsBF1T0xy1QF7q9jL2PBO0b47IZU1IYnYWrWUkyaso/Jy
2w1Uft+PAaxKdabEhhlqAtW3AIa1cHap3O/aAZ7Eh+BxTsI9yaRPvMlJ62q12R1qZk+TcvAnu4zG
Gdx1Pg8dmvRdORgtOOkdOub0luEE592z+b6Z4gxxqhY3QeJ8GSl7lF+gaVYa/eb/waCmjZlQx55g
lsAM6/lZzOvp0/viRw1sbjsQLBI9TX/3cG4kb+a71Y99l0Yex/Bs4MCx89MyjN0z56Nise6b0cqF
S8iPgreDB5gM0nl4JyXkNVJXHPymu5j9V2dOi7czE2sDCxc9/w7dIP6ghvy1+l4qufzTcY2EIbeF
57MCwAWVLY8ne8Ffi3OuxhZGujkUwf1H4lMUAoXLwkZcKIv4WhJWvGokVk0YN3MO/ot9/yx4Bbwy
djrMSZrC7gj6H/tUI/AveGlT1sLjd06BSSd+SYjXlAIKOY6ZgX8cgumj+RoE8FHYC59XJCPZvUVR
d4yuAWvZbcFeTdEczwnADXg57+t6KYP9RIxd4rwuqOz6GFty0rrEMBnfXX4PsBtVFpeEJ7a+F5B7
VE71DQHjOiZBDd2egqM3zDLUz1Iwxceth1yNjyHV9ecCtaNlPL58817RkYeAwxjokr3T0tln2Znd
SWi0RI0KFGk1zlqwz5zkVYsreXGhrv7Lhkhw6QPxriQ0jAaWCj1epSikmJt2L7kyA8btykqdfcFF
choy1/bcufzmDxJseBUS0H39ZMtaigCuylRCH+QV+KP3goKGMM1YNpcRi/WDhhrqzGb5uwzaJiMe
lN4KtDvHnjSvpZ4hJvDB0MKQrwIHRn+Id8/cZFIEGpaRsueVQYJyjE0OKSeJSTLiRPaL6WIjobxr
dc3Sod1zmuiIEv+4VK5lOwzCz/5OwPuCJ5miaqtOUIPDRv5o7FdAjmL6no5xYtJ3aYKTWRsDPCLS
NxA0snmIkdi2y2QEVdz6ihWp3wYEsWC1NOFlCezZvK3wEET0UX7nLr5a7aPfaJGlfFiHLtP+moSo
ceo12A+BnVoLw6wD/IZAdnVtZOaAI50nNHoq7dvkOxq/XTosXds3URzaYXEgTzBOoiQhnWGnqVQP
2fXQ1vSSXZnMdeeyhdpIT8k4tSAImtRuHdRmAWWYxwU/VeG5e2U0Pjc2rrnGTwiiPJMStrwbU8dK
R5X3CeKybhaiteVal7vD1gdFzH83I7qqubazsfYNfgvUFNyM0aXw561BoyOoY+8dZD8otmJgC5W6
D3VlIwpbFcd/3BgZJ4wcvzFpwEDKDPzASNZXcJPd1ljysHYkitzH7Nq8HHthhfpOWFxqT16ZnZw6
akr5EOCsHnPwK/b/OM+LnU0eLcZGZk7/5ZfdwegsJDFaX+6CZbRv8ew3iG2FBZi2iYyRqLpcp1UZ
TBdi9zBAIwsqOdRciS0S5aTmvA1Tr8ickfmgy4gQAU8MP2LW2AlLy5IaPqnspOCWOwS2u3Jn5i5p
tx9EEHBagvbH28KeOF66uk4oasoVctkfjOXUuxTk3do31VLIzgBmettiXC3AEgGsxK3MJLI5fFHJ
lZKEplCDuyp8KsJqgMAt/M6j+uqjiL1avEHB/wzA0RWlg6uHmia0ZmW9CMB23z4dm//3+/Q98N33
4aMDXkm7rTXYin4D+f1y90MowNp2fDTxJ4mu5D8rHBebseNVJoK3y65LqaPc0XUwIjmcO4oOdHjL
MFagcw1fEpmE8o06qrshuKjAH47RkcaG5ff2sWDrcy8iSTPDsGPkIuhqr4OnjRnJOk3OM1OYodVs
IP1jy29GaBGPMt+oS7RrBTc47fiPmJRsDMtlzpMm/kOpIbdzuSxw2dQMnoRHRhCL9Kp+8lpNYmpl
MlZ1zInzQdJ7dH+0+P3H1nDKHG0h/LP16aMfLH1MkRX9kqj7qPLjaNwbuCJsx4VxFOPdkHJPDd45
QZEEGX5dWHzqdcdoq/R9i9I34lurPdkn+TDS2992nAXpzzN+GnNOHaDooEKx3bXSdQNpSyiytQsO
vu1zvE5tsi5+GPPP5AOx7AxYHGwIZsUL/WwbJilKgX8AWWTm7hcggkX9axpeLQSS+kD/lkZFZdf2
atORJgceBUTfDGPkYFWLNh1JNKRJmZB5fZh7lx3hc0QeVPFt/bo+S5nRoA4MJgstejlB21gi3DAt
SfDQb/Bt1sZ9xgPDkC6o1Vf1bHZnY0Tw1wuA1XzCbOaK1lcSLlb/+BvUZd7N/iQReVikIR7bsbn4
7QS50z+YERIP8MF7fz0qgXEOXJEKcr0OhHF8kLDxEie2Uk6meZijyxaM/JBnKJLmLJIJzx6ZAL71
Rm7boCGqU/hV0WvPGiThTZdRHRp6xKOCoemV81HxZEvJMgAYH9HXHs48wPwMTo4KOf1QxktTdyXt
+mq7RDC9g2QoNJ81ndnuRIogaQ+e8V1dKg9DIwneZFh2d1LhTsA/JPS010I/evoWdONnMxvdZw52
aun+tnzE4HI4//4gMeaTrfcDFHbUaSCESQYlCv0cbhtADzwxV8wDw7JIbfCPg6UOJBTEAVsN9/ZK
AWtlE964kPIe8yecmfU7CYJu/8ItDC8Pvct3lP/IAnSHBH3ii+WTOmHhvIyxjxg3LF5mcUAafi9Y
kzMgAMbPnqSnUhQDaJH93AbXP64lrceaojcwjJep5rn4DvGCpXbSk0DzMefdVEToE6ejDfov9Cxj
lDcsbJYNcoHvhnSEhSTRNFgIfiCtRLcBb9MNTFTsXRGWTmskQppj7qs5Vu620VGI2LEiFykYsqNW
FgZWV1xuPAHNRa4LFpmjIcxVPCvh8cJF7I6FSoB7IXxbYC3jr+xs+fQ3Q3PsTBoYd9GJWA7LMZJB
/YxlLw2dR695l/HI7GUSN8fb4DSQ3B5EGhPlMKCYnqkMu278ytTqBFUupKaUz9Ifzx41EAzdrX86
rQfppH+zDqEfd2v+DmVw+qqCCuetNHUMwG80n9q/kUkxJfO0iBNzkgN3adR4Nwtr26s9biZ585+H
vBexDAa9J+PzVA+wWSYjOkX0CD4wO/wi5OGV3tFdOubmvb5HNeRvHH4JTFSdrCGkpJNxpJfk5Lv7
qqx+4spy+OK2XBSqNFR4PFV7Ke2oYznDzhm5eLtICgsMX2N4z1fQP8mg7+LA684XnjuEUDj7Lxqj
c5psZhEkg/6d0fn9yzkxJnKNsZKMQ0kt5KQWr6TsfxjBh3I3xgM+8282ACz16uxy8xGSnICo7EF/
dUoxeCkCIA8Hg+KeBHMC/K2+YxGn9vlHXD0dDVEABxwpLrXU05oeoB65g6MD9YnhsJLZ6440U2XL
YucjeKCg50dZOk/QPgN3y/KNXKDfHsJvfyXCpJkVON3mq3TaicE91POUbrOx3cwS+VI/Ep2Qrgds
djQqsXzQ0+HyUAm5Jec5weSP6BIntZMK/bVKmTgI0GZf/rIGrmAgxoAXb9hD0hzN1HgYLea9wtJD
pKd4aghVw4fg1/qiJwdhYPq/5UX6DgsQJ29zwR+bSo406ikgteLkgS2exXxHO6uNQSanAvO1cPW5
JsdV31O8VY6RoNumeaS0smSG3+UG7DS4QQcWDiozMH+94tz8lgfmKiZAXHdNFeyLhx1ayr69CxCB
1JeFm/nTcnsINK9E8axeZnbkip9btHO//g0c0dJNPFIPwyrI9QgqCAhwDY+7lhtpfw5TNadfYfku
9Psv05qL0/qSZFxBEUTFPRANkfu2Lw76VXnHos+yO/KROOMHor7bHpbHC6ZD6vvJ62a7mLvTWpLU
+z6z+X0AEseb819qB9yiHTRBWEDxR16upIg7KtVRTOJohIDD/LqEM5aRERQsvxqzqkaz/IEgY+Xj
eQAyddqJUygJAwLhycET4VRVMYgSG/AWIM98/dKIU3C37Kzb0mwZrzQUlfUBdE50tjc2BPjNnQIk
Kg4auSe3SE3M2F27WJH0UgjBUOFveBX/tTW54yGt/bDddDVfuE3r3xQ3oaF77AallIZIJKS9ACxD
a4l813QVNZxTEisu9ptUlXUPJpLlxh/JH7lCpR/luSuJm064B0VphpkqAmwbMPstPEGcq1qiOl6H
scyl7ORW+ovGIuUaCtsmLkf7Uzx0nl5K0AN+QjNAWMe0VG0b373TW1k3C9jT/kWMUDS7dWAou7nO
G5wxgRbX5S4g1nEX66bxZGR8aGx7Nq7wCfO86wzL+ZbAD6j3XzNxhyCxjQ3TPQPSKi2sgO9ya9Bk
nA519814TAda+kEEXg7ukBDRyU0KB3we05dILQX82czLbMhGBDiiOsdVLFjkT8ecat0sUPR+UZIM
paWnwDVL1nkhXpE7K4yUQ6gktmhrATK8j+ncDfSmXooczMdPs+SLtFZGOyozztNgCBoQNcbB8AhR
pjRnIlCZdy6IvZKcbn7sIt3l4/tiPPUkatO2s6QTX/Z29VyRMGDPYPQ8LWATZ8DQk3D90T3RjSS7
bm6ZU5SbQhwDSpFeD0p/6paSH1tiBf6jJrAa3ASWLl8v9vv9oaZtPzYcedwgoXti0IfMfOPlP9J/
1InB8ewtsBvr9E1JVz9PHhPT2Dj30vr3fgDvR3c1oAt+xRerwKroim8tyinFzaADL8VkOBUAu8wB
ZIEPll6dF5BiuvVSEb6UgO/lj8dNdR5QIrzl+uiAgS9UgKDXpIoW2Bg2jFxjwSPeh4EOPJmdkG2l
7h0r9+opN9xS6OrxleMZYSW6bJ0YnSAp98uIfok1KJ7UaEjPdjZNDvpF20gNrPINkaEREKEPMJNx
60LmVOi/mK7G+gZnifKdeKyW7hPUKU+idt8WxuPd7ueMHuTBnVtrx6hhiQYNltkbt+p7oN8Ai5oK
vSFfJBp3vdSmH7PkyK6PFvbewa7kojou24pQW+XdJgGtAb062r/kt0iPfYunZYeb82NOujbBdN1S
n4lOfLVIWRmPnJt99CK/TRKdMTiPEW1yXxTbQ7W2TH2LIDPVtXnXv5AoM0kJLTG1QD0kN2mH5m5n
nix8pRdH9csadSyE13fdUSpHbz0H1PwAjSbMpgyTWOUjkhkZ41mRw5xboCGtqtrlH+DYf67iQJz3
EFVNKVGG9SUuvPumUAc9bGEIKSeCIF7U2q1h4fP/MP16XuY48tKDbTqi9J1M+JuMYzJsr2+AtBuG
eoSQKGducBXhms+KSkl+M0BSDkhC2UnT/rtV6Uha3s2ioBp4dTmfmNxsmgd35Xn4UFdiokPR52Ip
xTbIQFZcfKZD/BtGlqPTAXNq2gLiPmYAgNjnSv6sHHc5P8FTMXrxRnwzwxe1ASszKj55uuLo7QBT
iK5S3YHl/h+cTswdspqIEjvs/4c9L1xb06BNS3/YnzNGBtijjcfB7orKYG0YWmIzWee2jTItfC27
uhZMSQeYpOtOlWhG825S+eMuq5ZUlSDgcOUXqgQdXEnj/EtE1Shwo0OaG1j+KBdjfA3V+hyjc1CT
cp+lvsylbf6b+wuEVbZygHr5Juynp0RWELv8bb4KG4h5H47aibiSVAYwFW2SMZS2+RUnaYGTaFo2
tbGL5PRD1iVU+rgNCHvRuqUIr2vTFLANVL3DIfumDxROZ+kks3H/YzHMSZaFH5+vhohF5sqQsgcv
IYdismPun9DYJ+1OX7NDhp97j27CN+d1U41WVT8JXKaLCT1QXllAg1X4p4p657If43nblIEv70Ix
FeHj2JPxX9b0qmt0JiCWDJDLDXrLCoQFOKcMxlsmQbA5UzEMy7rFvEIjizItKuqohjcPfI6BSJBn
ZI3WS0R3rqnyfiAvxexKxbMhWJ8uTS0YwY37tc7suV0+vhH4TNGkDc+NvYD6zH0i51bOYb/QTc2X
Os8M35jeDGj7CcEKZEaJS6ogBy0QYtU1uGPwH9uVQinceR+uGgZD7Q2dgfxBpUbTpk0+VFY6CpBJ
M79dNAwrf/MlxnBTREAPwnQwXv/sRSqyLu0fXNJ+5WqgyHqoLaTuACZ9e9ygA8Iz0TTERRNwrXGL
lQbPHKo5jA6epSqLxcTnEBhPRIHja+Cy5jUucTCytZbIElvvBRRGlr3OiKeWyT6+5trBgeqH0O+B
rua3aPyzg85VHROwR+LmyevztFINTQ+nh42PZ4h54h+hnQZt7lPR9uTgOtSXN3d7ARvHFbBIdN4G
DZqdd7kQiktG4qbchOEl8g0CFIWAblqowWuvBN7NBB+pN7H9xGNbchHwIrHmYWH0N9ADjnsXn5zW
bFph7LtPoduJwN+Pgh4UcMLnYReHV7FntucKyqlEeEdvR05dv5lfs2xlURjMvytSsGyrKwBlnOht
BFQjim1jgEowF7tL8q/CWGe9YuvV47uQn003FgG4/Oro3ALzP7qJjGUIRfALIMRzzmniYRZF4zBs
Xd6XMsUxc/0KayIMeN90BmtC9ml8Sqn+2VkKbGFSIM6KbTh24Gu+rGbG2hZNEWmUjJFMbOxpB+pE
v9T2D+E860B0ut98PbrV89GygYFWXO+QRdktgAENW3ADkYxnEUvL5hfbbOAfZxjOOsB9yHfADHE/
iiFwR0nvoJ4vdOGdVhfRFUUMSpEYG1kXT3KJPnFVLzYr8q2nxDh18z8u0HwFuve8cdGi0Zye9SkO
hWL0c5xp3xH9Y1CseWhRRiQyE69wrlV9D4iW0440rEo9TTGrLSE2zYp/ZbidI3RA66zGQ5XfnpON
wOSxOpsXRkAMzVna9rRNcjzhn0+AXF+L2UzE9AibKcsAkQHP6r6Zi7H2mpsPoLh4/9pw+uun7hlF
FGBBjXNRlfy1ljzmyrBA3DSbVFxKqDHb2vz4UCKH6XUAywZCRSXJv/kj5UsB4PNdK+K+K7LAIvBD
EECTByksWVw3JxWzf4sRerXV8JfnXCZHkvp1zH2ASSvT2mLdtjFw9tfr0rv3YjLcn7pCZJeCmo8p
ldGfO36uOHONVg8NBW38g5DY3Dg45q/da9qHuI2QY0OC6fcCQo72H5IgRh2+LXdB5JZvWd7f+OyU
3q9/LlyuyhA64qUERZaH/3W2hyQOjaERs7HFuu4taptVBMNo0023CqDhpTU0af8oErJK5FtzvGTE
KkMTbOg/SK6/ss7L0GeKFa0D5xJY5WMIa0FSrh4O2AlNdDxrByFmwlMl0PrucLRvRtOno29ODH8T
HZIB0YNyA8ylb3t9+VIxw3DwonMci8TVsmKdeObM/cPFOBYH332z9DiLNrMQtXQ9LsXAc7gBMATK
6NGR1IooTiQ4ft/segle6+IPdpzFKvWvzXryEpGeVVzyfz5diwFlp9H/ZwcAKKcq2huvG0pNYpv6
TXZ5dLtJz4shdIN/qqr5HsrNhRIb5daLb8WchxFsm0nJMt+xz1yiHB38nVfS6e+RZ3hM2iZdRHCP
ylUygXCG/Z4tIA3FsCaJZjNpM3zXG0tCfpAcjvgUgcs4StJ0+9MBTSP4kvlKsMS9i1SXGNzzNgO9
1FhQwdbyCl9D8MCQPBlpo8pK/7lCXhTO9cqL+kJS86HOsI1bqYF/UqzsHnYrUwi2X1o1xVPjOywY
16c4Uy/3/VcgHIDmr0rdJwL1Cc47dW50CBz4p9WQrl71APT9WF+aSdUTLdENuhW8mUTKla8TiX7h
2kYqnRAju52SaCMVByKO+e0Ade/bmgaIioico9RXs5qVz+kmQeNQIGl355M+HsTsLXt79/SLlmyI
aC3eo/s2HIxj/t6jDukxiGkZO4QFb3DRdf8Q1ZT4Dh/rRgTZI3fJ2Relb+JakLX+mT8ICwcu5uRe
dAIorYItyEmrYsgIeh8iJkOg+Ya+DnjTTtWJRv2N+D2ExmcLbfGkmim2x6MoFNKX3jwA36Xx3Ped
8kXdvVolJvJQSkkjMm2gg7evJ7IKod/7MUJSnEq8MwBjfkbVNfH9jUA09bc72QM8pX+560gIFN3t
OTopZig9zQSQsYzqdLyvHs/Qb5zW1j6rWq4LU0VPSC7/mu7g4LnADqQLpiC128m79Q0Mq+WeQMd0
GQBMtjKm8b6YQrwonhLQG+Zbx76/jIwyWVh1tldUdj7Ogx7HxKrnzTF7WT/5Ty7knGvcMq3ciE95
mfFIIM0CMKVofggVDlcOk4vmd+JayIdpv1HFuJ2I1KTKRXe2xUquSUpsSzfS4RKNVczNNSPcbIuY
S2Yc11i0lS/bL6rbnlfJXhKOrB/uK/BbvLAl+7CR30cDTZ7+A/doZmsvHuO0QGOGOK9v/GFEQ1YN
Fyz2iQ6yvSRJIuTMk7t+jL2+mPeVROIVAoA0sIxplKNBHfKjkv9TmkbXCocfaEKSF3Fw+B+ZBknu
Ngnuc2DHa8xJzHrB2E+nmbs0Hkhp10dG4azOIJbI45GTy+pzBNhIZUCooK0ikda+FKTHqeTgdCHp
YlXjyGnwJy0e1acS9t3v1wCFa6PSaCYjgR1MiInG9vnfrrpAhrlTla12obUiEYLXPk64e1UM1eOE
4iBXBruR5lgWLTEmN+WePht06SXN2uU3qKvsdvM+RmrqIeIQWnyZTqLz/gMh2oKNNiZ6TaFO7k+3
TroGKt0jaJAdWBfCW3dIzpGpprwpsLQpUMU2UdNmgb/JazNSb7ibEc2iICK8CE5C8fBkB1Zcvyb2
Pof+u/Bh22uhLzX5LMQJ8gaiTOQgyTNOAVL9OyFg1GFTuKm+DZHGuno6XVnXzIC9eERgDUVx9jSi
onsO7b8tLVVOOvm8uktb3L37BewSbMj39OnuuHhs5gMv6gx2FarECvG9g/Juxhy6O5ju9CIeg3sA
xOkp+gSeCrplL4RzRTvkTkqaUacdvnUtbAuhF0j3lkBCwEHnPXZ1SSaHgxY+iA7WNCFOpxlud2Pz
6p04OqfAMX82q4UVfl9N4iLQo9+rqVaI3B1xkWABvUml52KtIDlic0MHuKbLWmjJ2AV/nlaZfnwB
Nh0uYH89rihsqPA1hMajHRWT6ACkVecIxZt7AyXSN6jEQ9j4rwcZu7aRPRKt2MoyxS56WqP+KEew
lA+UCJMRr82y3wRLYCJ9mklbLIyiKyXbKr48h9s8UVb/358Epql8lLjX1FFcJIS7cku70bFddnvC
7bS1Tx3wahAy6Iy9+hZ1Jl9gDWRtaYVfVNXOMRuUhZM7/l3LskFVRqocXyv6JMLuQzMrLNKyAuSd
uD9QPxjCiEXbiZPYGBBgiiZ3fHTTC74A22ze1ZbAtVMKe+StZQy1Qdiaew+yLzx2/J4oo6kJpt5+
G6O0nmBGXGk74AY3Z+SEozU3Aibgzij5ZXQxqI4vOo8YaLZ5splkbtMD+uBl58usApaicD032KqS
Dop4pGxUg1MclBgvSldBGN25Mqvobdkd3/cX3h9N6aGlJnAhpww92b/NvGCsv5NEey87i+HC6yKu
Ds0kEG0/8ZEr4Oc8evMxuujid9fCvE1nJ6vQVlVUFikvPIvii0TxtUbjktsUBQ/EvRnQkUGY9Zma
EUtwHKInRQ1A0zzjuPprv8d79LwWK1sg9p/Qv7+DdWOAiLRWWFLdNPr1Hhne2W4CGsIncBScglCN
TrHCpY2mnmFCxPxbzOKq2olLI2zxFg84X0VcUCcY1wUug8HtkLFGwyRk52+1VX0CDKZgn7g8T0qh
53ePk/JaL4qPIa4K+xgCUslMxb/EhkZV9iEwZEb+WcOaEhtO2JrrgTHg5+aFOCFNwAvuFRjVj8eY
vovLYgY0+r3y9f69Z39xGiUf5TE8ig+1NU0VNpZj12ki5VjTHHe8AD9wmVsIdWw8bVEqIkrM1eV6
nmluoOCBp3RBBrwgtXnXjgJxPy0LKceWdrDqDsbukqPrULRZhESDZzXRcyw7JT5QE/1LtQKidAg+
kT/pYB3J3HNcWGaiep0XYUcbyxu29k613vBbIc4lyTcf1oW7qGz8XBkEslGXx6bxk0D/CcdIRhr7
Xx+/0ETf+hwdpn5fL5yVDIqBAiwDXUfN70PCZ3BbRqipmOPqqUSL335HgiVrGLOnEW3e9YI9bjns
3GzzxSpgfod5Pu87M9WC3Ghs8/MUBy/ZFAVm9fAQdqxAW7L8knrhBSckt8Ktqho6iGJ/+ImZtC+W
CpXCR0jHQozL+OSqZKJkBizcl5i6k3KX2uTQbkE+B4DzVOyVTmM6ZmMhMdwD8dm6YdfrGtIcXn0t
WGKN7HzUl+c4zmDzvWYg6xXV08DzMGEo00GfKx5QOZ+vV8XbXIp/9eP4MtN1nC6X5GdYjnQhlwar
Nkt5S1LgYpAgncgbScsCW4ztFeNI9iDIYbDJ+32v+KbqTD/f7/TgcH+qAgnIeDjT9S8JjHVOJM3I
S7Q0ZSw0drAe24cSivqknYLtr9USBBFcblPgR4gnIO1aXnTX56V/v/Pqv3ORGEMWI65jGimY9xZ3
vsHjqIEsiK7Kq/T6uail1S/slIdefaqV9702EPufIqdjWYQhbAivsIZfj4JiaYo5eTv9IDjCJZ3d
hbW+yhTsFSH2uZxwQfaepXDJ3kw2m6Doi821XXAgEQ6HgNBVov/8y0OD8xq3SFRJkY2vMglSt0nz
FgmmIiEvBb/Yp6nOOLu96p6dkcuNBcRXpnfU0IYCpC7vIeFN3gCeKHxDCFaLzjX2kmz6mVVFNlw7
Pge5CdLRw7hivr1rTtZ+w/ICTzeOhjaS+qukihGw0CcaxQCJdaau/3z0ZMAl3IYs1RqgVHXHFJKF
/5O0e6d4IxLNFu8C0quEvnYk31wR0BcjOxSkZ7GuEMkM2UtWOcpdVUGxQ2zo4g9XX0zLZO1R7EtR
EWz8N+w6TtXhVE4FPViPB6irJLKR2+kap8U0bRv9CtwzUTumn9v4hcGbeNG07RquNWrdJDBvWNOu
tOuJfYCs5prg4tmOoadO3OnLJYwfJabiFshs1sXAaOaQnHXtiGdd2auk20qeRR/ENXshsh4mXuJJ
fyUiTWdsw/IlCon/uIP+VIflgr39C9nodVxeAmJPA3Q85Kp/Y/lJVZV/P2Y1c8yacMhI83C1OGOj
6WGwCswNKrjEyFMXH9jbS0QF3Z8cMnUkq43c+HI2Ys3lr/PMByIhJz7LCz+BWtpj/hjLJn/OjwJF
aVcnAuTfM8rfuWr1djO95bW5+A7TQd3qh+Eb4UoPFQiBJ//xk1khJePTzRuZ8ps8Q+gFrAtKwby/
TTV2kGe6UUuV6CHwTTVYomrKCkVJbzd2Vug7wj/swA7pncFPS13GosXPAFoPV6D73kLPc/FSG6Kp
sqHJ7l4FajNghTEe0tRpQ2NsZXHxGS/WOz++Z8o2E/Uiwy2PyKmCiq/pheR58WlnMYSjPQBb8nqP
3drj91DUVR0moXvibh8oAbI+yL0ISK/P9656Hwd3vtxPV/WsAPQjF7gplVQLNSXcn/5eb+7mp6Vo
rJOfxPbBvNcep+tRnGyrOJvGBlLd/0U4OVphofAzlz6PKacf+7TXb1CvdRj2wTHZAhUhNiVRK3ry
2TyqlGHwQDm15up3PoigyIFq7/uJSMkdTTfiqvy7kVvqx7XhuZQVOOZ4h4VVZHlZsrBbrRdjxTRh
VgJYT0UVduo/VR+yzMX9kzViqFue53b4IY42TMo5hnSJr5k3DP1I4f0NG7G4SABOZGRu/tNvpMBR
eq1hQvOJ1mG53TXcZvkbraCK/jxKj6GKWWw7R9iGqCx+73Jl1CDkePd3J7k0mPUb7X4/2o9eF0Es
RZ8exOCrEZIWC8eNzk+5fJLYpLN5eJivVFW3FeoXp0uE2ojWi1Auz1ZK0cF+lUIgUkq/ESzsbM0X
Ige1gkue6tWtrsJVfabkF8oiHtcHsEtHifiS7oiuSRCoVwKas7UbR9Ov/TN5H4H6rmHQNkCN0jeM
dS7Mx8JokA9fv82nMzxGWOpUJ8yRSo3KP4LNP8TPhZLooRUfRETHaNRHss1D6WxcB5IDlBy7llZ0
ACWy+hLkk4incNZA/L3Z208lgjf43Z+/KB79xJ4wko5IOGWPbyXQLCJpEX6AXyB7WbfbdiJqVVuN
bkKdUo/p5no1ijbSh+fSEDHEik+twPHXCOJY5PgSrPIrtgYmkUNCWi5TduUks1/npSNrLcD/f4bh
RSgaqpkfjSLt37fwcJ4R+h7hsuHaRSvEi0lLv9d7nqmECVVyRUrHzFaOG+c2O+4x7Iss9YLzQIAg
c4Mlr+w2LBaN3TX4Gw9Y/jTcFyRFQp318xvPmxxJdWm7/eBouIbqHCCVemiwA9boopvWvqBjctCX
0btT+UG1xQmbSaeEi7NS2mC8benI4aWRHoy0wXpRGgKhWAJaLEB0HlPjQaeTjBDZfXHYFudxdG/x
RVcrs/xPwEhheEWFTFFddG8/mozNdF66p6ZimJZNRk8jgyyF5Bi7rhNmWTl9pjd6IzjUFa7e++Bn
H1s7c27iqdyoaa0GmsQYSm/vXQe2z4oETvyemcpyMUkwX52U1wMsruPheiT9J56dqizLuCNYYpYc
fNhoRj0Z/aVL+jABa80652wPleOlYGDWP3sOqNQL5rZdgacnaPEoAwrrGodmwsoYeExvnOQP/T53
Te5n58ARoBHRMjopFiK3bZb1cWRpfWrEv8nUW6dgm55YBixrITEii3hDMhPovo36j4DAmhE1WNCs
dvVA8ija1vx9djzHQLdkemEt5Vk9r25In2JlzfxXYI2McsyjaMTAIT+uTgZBK/AT52ubQeANAk+Z
h05pa67kCLcXVj9Fh/NdWBpgImjnjClZxTNN/vJ1p+CRQXQdk56tFiacKjaYHrURLZgQ2VZ2eKAf
v0fMW63/GV930TKJYPVZX1zKHLTkx/A5wAESB8ow2mChtj7dslGl4ExPeA5ZrPTQsvJ64opLusM5
0sczBMSo49NRoSjrxv8PY3QedAxaIXt/6WyH1GGCkTn5QC0MMo+TKvsR0MdS5n8BR8s5HNRPrUQR
zNznJVaLoKFoBudonT/1b1JF7SNeMX+DOW7uJaQXgW2jvot5oN+1b5xjp0J1gXyEE0HCq37Ct85u
bQKHwMYOKVMWQb4PX5hfQiY6jN4SOci4C5RcuCwtG/ZZ3H8Nw0QpsODQTThVP0HxZkWJkn88lc50
K6wfkIrZ7Hj06Mth/s55FkPDsluYIZJPB7q7IjuALCP7vbI0ruZAyTZWDbE9U2YITFcVnH19Efzo
6tB47ROlt8KsNpCVx47NOMY5xvvVW7dbWzGtRLAbNmd0K2iNlFaVaE23sbVCmQjbOLMXxPDVnlQN
mFsqtbOvkpIMlg7bNGdkOicF5voxn757LFaUSdl2SLyA1dE7RuF73HSkBrci/6wbCZgGXGHafJWn
T7ZRcwluvQG9ayxzDJ5XXvTZcU9jC9OL2HzFRdie1/yMihMeiMcN2zIRe7/2uWOiU4JOvDMPZt1j
KkJtPEvftaSfxuoXEzr5pMpQ2jL1i7EXjjDKLMl3IGoa92D3evFPvLXIpFR0o4Q+tzo7mYnaYsiW
qGng6174UFzNbrwNcbAXCncoWd2nAed6osONiDGxFpMX0JjLP0Uj00wBCqbGRGtKRorxMKTGGAup
7HWzFBeZUIU0z1KNvAZno8A+E56YOlMm/v+AjfrlO9uVwVv8Yhte3NBeIYsTQJoJxvBAq9IxEkIq
p0pfV5M2lqVRFGQD6O8IL8txPd2S86lnuXLdCc//G0+LB6g7Tm0IDPSgoc/ThriJy0OvEWU29kLY
Ti7xpgBJjF+Jhgcf9TupnbcTKeJqtMs4ijnfjmgfUYPB3eVtWlxecUFTvFEiG3iJxXbBXoUsT61/
GreS+4F4g5D4DfwWW32G1lk7gqr5GuZzU09PsHclN+4qEaZzVqMggUyoQ7pBMR3Q1riRO1D+kANU
DCJ0VoARBFmOWxOYuP2q5pwHtsaRdPkJg4IlVVmprfUgK6fvoUQVInK1AihmW3R0NGv2RkE9pYYX
tQy9bvEbQWG9OFJSLiFUxmh8qp6Zf4UE//HkcYZRJw2G+BnOO66v6gbwzDOlORsZhXOwqKkYVOg7
IwPr7wZwZxvIJia1Hdxd0o8A+CKmJ/aq/l40NCx5Ydohqd8FstYTkclWgFfG2iCtP3nwpBSjwHPD
osxwkBmANbTjEb2n+p4lkvUJHka8zMv9Z1+72td6Y3k4/XTSUZBU3D6Qa8P2jv4B2e6edqkDbmIH
fT6gFD3vwsO51MJRAGC7m9liYhQWZaj+lpO9dkOVK6ZtBleRxu+nvslEjR3rnwP9pCUhmB8Pa1lc
Z49vBc2zpl+NqIjDZSdMlxhzQuigz9MncuIwHy61Ttfe0vnEwPuizQWTs6S5iesjCDmK2x4RSQNF
J1Is82yfLoiVeiDJOWJKCuDfKCOZCEogxh/o0tgXgbCh1+A6V1RbnAiXPrG0x4cYsimhbXcQTa0U
JA739IbUYNDs0fGrQ6fdb8QQEhSkxUFthoena3o/t0W2uvvUuDuVGpEFapaysKDMRHK8dXrkdztR
YAmFnRK4DH1limX14kdQ3lX9Yhaa9C3AgWovxyvUFcQSJEE+ERNrTtC+MqA9vjWeOIKcHFhu8E6o
0C1/dCE9NCwZh4cZDnMejXWDLPIOy1F5T65Mfwq8+ZWGtzRybVtl9+etBkwqiL4IBc6JpGwGIlfF
ddQ7CwGMXSgqDXpvGgLYLb0nRMQ1b1pLPE51/D5heTeqdT11fOFU6811WdQC6TyipnHN0Jo3dcJ7
bTlubt0bdD4t4g+6OfjI3s2Xhg+gpxb2tkDkgYY4pmUqiO4+jDqRa6ztYXIrVHcb+BpZFW2+F6DV
1ybhL4q94itEpLIDpQNL7pmz0E2TsLeLB90HuNmisKXmw9oCGVVf0XRPzRc/TbqmgLFr4ZzgeJ9i
t6qrpDjlUaRNk2QHKdMrSeSShCSbKVkPTRp2bywyEIX9vuzkQLO6DgXd6HMjQ56G1gm820JwFAbW
vvABXtqlwFDnQKfvgaEwXPWHktnMQ9SLBWTOYLY4mGcNoYAgJ4hTJ34jMvITr4tocngCPLAurA7/
E9Pbyua3RQ9azemaUP5Yi09V+g1OPUTgkuSxglhpFHN7Zc9iuIO5JI9favNejwNcK61aSSQydXQp
Dm3th0atdjQrKC6vTPjhnJKLj6+CGAhAKuCAGgBKJUdqi5eZXBV0cO0DVyTN3O61u3g/RzdAWbap
OkmBroQ3Z07hUCNNwdXvnqdVG4UwzSmBnEv8v7nlaqsNqG8Ysidhi5quyA5yO6iBTexmvw9UFmdg
bFCIWNuShTDgxEx/iW92/23SyT7mgm98221hZX9BtmfPEs/vjYelDH006C15k41Hlcs1v5bc1wGs
n+GlP90Bil/HYYaHwI14w8sNv+AEsGgUdcNJCQFMFZViqIz0ApTQ1H6HrcYZLOgznmxgPEVJKT0D
13R9RhZXbP2yfzGgUqA2D/zkbEF2jKprI1COGQI8Ew/KJdd+UUAZ0s6/wB2y041kbWt3ADUBiRuS
iaMIFCJ7EgFb7d/RyIaZuyGcNSImte4EihbfyXL/6rpPzPeRDE52ZK1F5BqfJbFo5JlJRQeSI5+O
5/NGW3X2DYHiIUEFSlOTUkI034+xcGAtL2Kzl6bkF3bsQHHM0GcsBm7JG4JUd1fdpu9I4oFkDhK/
H+DGpfcYVDgVlsBVn/RPlzePIv9l118JjesM+XMOhuKvoTw15ughjhiH+RRLXSzsSBhMYo4uBUvD
MSfzUX/WRvz1kWy2H+uJtpjbjQkws7Qf1t9GPdVe2iyoCXE0IkRdAOh36FPPNHyzAEURYZYnXp97
Md8R2OQZZ888P5nsUgt4aA7GPGN9NuLyzhVKJv3qhgJf9uqRVYGSzVT1/GmKcFjHTY1xAKkBXA62
Gxx3SBwoodkZXo0hDFgfuQiITH2hJr5K5r35hcAPMNDFUVUqDIJsEFC+PTybrFmHf2M4eMoQ2WoV
5B0pCG46e0FLLRVzMd6sEp/RYTNV756lc6oDYWQq1y75DPmFA20Etm72U0DiExCeRBbbyX1+GLnW
wQY06b1ibz+Bl+EVyv7ZENbDUUj5lMS5T5P9Vvz43nNt7ruMXwjRww/8Kv8C2AeckQ7NDm7vRRBM
LrxSMmpuWdi3kIOxax/p5w/DUhhkO7YTSGNPlszmxkb89BCWMw8t/2lhJ04Q8YPtN8zqNWjkn5LM
J1h14g20Pdlbq7WeqE7JhuQ2BzCWvx+o6svYop36TBdkkBnAKFdgGMnnnHRUZhxy/fLwq7N/8HAB
rpzpVcp8d1yHHZGX78gDXyMel4nYfnVt21vxEJPXx0io5SZV7cC+9lSeZsw5gkbL9B0nSa4hM0i/
CQgfD9ZFanWiXkRVe4e2GptoBHSBMLM+zphDQChIkUf2IC6JmWbOc0qzWu5/V1uAsOMvRPljdPFB
UscihxwW+kO3Ik1lwePMQ2wRWNR+qe8cEVZSLNT+nvbhmaBB5e/ghDvRJVeI/EOx/owVMOMXDLw5
TK/B+LSNGaKhm/PjUOoFH8TJ9OEFOXgOSC/F7DJ8fsiDZFBWV50ajtVBkhhcajMITB1ljawEJjFf
Nsn+mWgs2kfFyNaZvdDylbzpbPyXYAUceIYIuwcD7Vu47XKJSlB+3WtoDDb7wlpORy3+ekB1fEDY
GiU79tpwe3n2luz6BVXaesQogf/Cg07W5eDb1Xu1abII6AHUEwKAzEhf2N77lUyGsB6ZKJg+1P/j
HU/nxep/jh9/pstBORqmsSRL9lGrCRBPd3Wb0IqIAUvjybk4kdy5iHRhczWZQ3CoU6IPEq3FllaE
LuKVS2Y20Rk+cH2sFZN0paJe3vQYJJwl6H15SVF1v7VdREvniBR+oLlYaXeLLDt/NV3qqwyL4hf3
mbDeln3r+aAo4ukU67MjWJmjv0zbsAZFZ9gLK5b97mv5+UiNWRQE6i7tS1Z1VnFDq8mw69Bf5Nmt
eh8EBSdR1+UdebMKh/bKNTZG+h+1K90bLm1F3UddBGgk822sAi4X7Z9JT8gVFmQcbpmwT2J9meF3
KUqFKX1lfsgWdiGPMwhBqvn+M4VfBJcmxZV9czeGGjR9U517HEELfbTG5Wql4Xv/E+3TlTkKQOoc
3+x94206kgWyWpXnPJ11hAmmxBaqoA5n39icGF5oesywr1buNiJZ+6112IxIVzBgky9r5YRvU72D
VKNHOVQadY3xn2Lgi8ySlgiiR2GEyBjbddGZTwCcqMtYQBq/FXc7wo1KtmVG4gOFxqgbxEvnptGB
d3tOGkXeHt5eL0qnVxJ5HIP6mLGqddzor5llF6jMeOwbp46clLcX8fGc7E6WQtigR1dyPJoq3JC5
N7RfWI40rLaUwOms3E+QzvtJ11jVCEttS6DqgnWtlpYvLCtzZvecOrRLJm6VzTCTIEQUyoCs1Sla
rqrCi4UfpDHhGIYGOx80+lPRj/tchRCGfwPUFDH/nvo+4MhseWeYsaPqIXhD6rlRfzkw/alp1/GH
G7njTcxJBhUWGCzj9pZOSW6uEIcYMGopXs4KTnss3cJtttiuttbWSZbvI+TJMXJCTLWZHEJIdHoM
6u3M0+SHm1vPcP4E7zDtkZeQSQ9JrNTiEIS2nQu7cjHiP/NamFYD1XlIPRjU5rl8T050MGMPajuc
pC8a9ZPqhvFguDcl+mZFavEZlfltz7Wm6zppHtlHwmxM4oKv8AGB8ZSgMEgYbkjGznNVjFUkmvoV
xbl2qFc4m+5BZIl8OvusTzjS4l6Q5KXJesBMG3FUrKuVakSlc18hQrLXWh0Pee1Q8NLbePIRicOS
o20jqzG56Z12ag5oyxR8d8HTm344HOSVUiToo5YP2JnFfOfE5VNtub4ZlhJ2gKWvhx4VQhHjPELh
jFCj11XEvhz9aMgCdLwA5xSqNDytMKE1vHRJww0SxlXpbClbt0V7NlZ7xrtSIMdUN+6F6H1Br0fu
h4R+HhRtSC/eXd7BCwAtO+bSCDV6iP/L1e8DXvVacaYdFc1UjNjhk7Zs5eiZ2P0syLY3b1PHXc0i
49DIjEdLOTs8ifZA0a0TFmyYOmAvHyMKXWkMnGZU7LuVPkjSO0+zHyLn7dMuq9+MqllTQVaRPMvZ
pDE1Zly5xx282C5WXkyskX2LiUHjXjVyzhiXG9MviWk5mRw5QcD9AeJc6btyf5YVj15Yd3oazwwr
wMOb1lPTsUJzjaXHvTTmPEYh2U1uJviFgEbHWt8+XRkOraRP65u59sIvmzTGq//L2KxyWpNku7ZH
PlGTEZdO/5sa1aGtnpw2cxdVMA4EzcvIW4fh/AZiT7TxyTyL12ATkWPkJQ8HqmjvF0yUHeqsRgYu
6Eqb/UJxHlU0xUmQ5wUWx8IOIuwobPC0aN4fgFolCO8OKnkYfm4DAYs7hlnaz3//5MEzax5cwW7O
odAEMc15BylUEtG/va8160JAOy8FOBfVoacjR2jXFjw+k/eJBeedRbURswDJ34+EUZC0YAYhOQUL
o2SFnJtE7+glin45+2+oWbCmwrsYOu4IbfQjl0NZmS8sA4AWGd7IGq4sgd9YzGRZ5nG74rlOwAgx
ViSCkNO9AVdyYogZnk8PWcB6+kzXVGu+bm9vyKuMGsjXlCsvBGBodhQsiSuetwVsx8S3GC+v8Hom
e7dYjh7dp9xvgTcXiZ5R2PIhOD0/3o6uBVocaFFMKix+oohky1DTnpAdjjAh4hA25o9v0ACQPm5/
IpetkaA3x/mHzxPeeGSCFU65TR7GpIDOrKb5p3TfQws3snR/NgJ0nRHYcg2ZEyLVfNJeKjukMGFV
Dr/MJ7onqgXCIdfO7h9rstkFOTjUzkBgB8yRXmSWjJ4m+4+J2OI2EJCDXRbVrmajAFISWsml/i2y
C2489I0JIRqGzyBuoI1XosvgoNYe6bbKC7ZxXpq53jukF67pVxjC+pPdfLcJ30SB3TE1a+Yw+ok7
s+p7f9xR8LpKaAHtXGqCV/l4srYb7/x31bNnT0VvTqHdLlSA3qUP0RLi39UZdAA+rFQty1tdj6Ld
fDpOGaWrsyu0fdYB+gtmUcFm4Mtr5n80r+Pvebc0TNnyc6BH5smyVW7UJA8mGYMTw3kxRpyEQm+Z
j6Sii5FdBuE3sx7HGxO1hYYx07oSegkVN8SsSD0bH84xY+tSlhSf0Si6im37AtMEviZpwgWR3VWZ
KG8Y/6oKezXjqwQOGdd/YDkOfP6/RVxfZYgEB/yK0Gj1z90sebHf4+jqRzaPWaaBT36RKOncPAuV
gJdleXlXheerN/81jiJ4Y//qx/p4Ygvwm6brf9PVa+FwQ7JnGq0aF715WVX9W6gVrUi+8Skr+Sdy
cer8gHqj1x9TySAnv+azp2ekKvnZR+xFngC0lKml42pnC6o4CTdb3ZMaElws6zW80/9I98J3gT7u
9EHN3LNx27XD2v7HdYU/vYSxLm/CCug/xKVyoaNGg5iXJlL6TRHpQBuL+GF6HMIGLmGEx2J6lvl1
ZoVj5VIM8noKu2tZAfY6vIbXLlcH4ZJsCWXO8JNWMwLZdZL50U6kLtc5JnEgvRF8gMU4LikfAlBj
GtE7zZnfWS2PaiMZin5rdVNMbP+tCUM/oqeUXwonsr2fAx71+8MEnwDXxqYCdvl50OMSLbgdCvJ7
EAzIUzKQgToWXHPKrrTYKo39lNSQSAPBhzYkYNv7GCcBSO0UBQRmcnlGsAwtU6EyiZRfCXplGZ1c
qJ6GDL9ytDsqLX2cHuihRKUmvPyu4gVz8rOXDK0YR16zrOU48CzMuBgWVMexQc+wlzxqlYnNcVFp
b/z4sZ27C5upKB0S8AoalbyTyE+4V39wTPZqrPxA8C4JWPmkCn99A6ZVRBjgtKuFhf7FhnygSq+L
3n7hDuOA4E8Fsw6pECBgGbpGHmclRbnklqH/erBtO2OoyFKFeXRpJv+NeKjQsaTQzfoiug/Bs8xn
rcN8WZrwgXBGTtoBaiSmBtoW8FvN7m/9DYRhTeO8x0jZEODu8EZ6I/yVHcDBj3VKj2YpFAVjCaGr
T0JfT4n7Rw1k9xB2xgAeETvklZegq4lkXusvkP09PGP78khqJQ4Zf22kSqqfr9JFuiwlthmC8wg/
f13SiIQvHTztwRNO4hXGFkkphUuGR8SSFuPbthpPJJV0mi7feuTFBh0+dANmnaSAibvcnVuvnik7
5f+39sMz92jap4+nrABl9THKwI7U5YtMB45Udn5zr9l5R3ozaF2uvHIZ3/02rTpPG38lg025UDFS
s8SLC/K+L0bwftc3xz9enDZR+NxogCIAIK4i+J6nZ2K+a4X/dKceMdO9ycVwzQG0yDqqt7TfRgBH
Y1lu4zv2LNRfDNp9WJtrdyLpE6VmeExS083kccsC0sxbX0873URVxmH5jBsEGttg1bO7lkjddtux
pG9QZwsDA1x7YqD5/KMsCFr/WHJ/xUG19RKkauApsITzuWhPlDp6AHBx7bhmf3yLYx5Vc4lBx+48
3s4jZVMCZBwzNl1AocTELGTS6o6T3fIKBarZGEkepaYwj+T3OWQBHGARF3Zu621aFD+W5YCBWYKs
aPwC3QWFBuONCu0YL1CVpkKz7/CNaS6dJINDmkbgNT3TPEjwfdNT5Yi4DtGsmnOqvbIO5RhFnqQS
c7VkIOkgib0fmwSKBZLGhdqBzrs0X659j8vp/RgPkGgZtjcutu3klwdBIcSM/BNP3T8RYlX5eQkN
gUb6IHFFqpFAyGDuWAy3m3fnE1xaC0lZqUgbgu8FZTJ1+opB+octLPSssmWrU70JnsoTfQAw8848
pRJaV4AGce0OM23rHBKkpNkBleTqldSFbOtTsJ8bvMubbgOn0XZQxf/5COa8cus0t9dF8IPCFpO0
M6Z9lwQCUwWFpgAKn2sb/Xn8F383//7GlAtHBbeNSEPyskHlDmQ19EtoDSr1yk5sXOaSF+dL+MzK
fPjKgB7eEptOp/Du1+vPYMn2aj7eGnT1Vtw/YpMAooYDGxlJqQRqX1fVBLdt79hOkvqjAnGqCKvi
W33NupNVSE2Nt1KVGh8Cnr83xEeytr56Im23jmEBK72lV5nUuCEnCu8JfJLatYmUdR193gFmsds1
5CmXNY1ab3vpEISSNPKgP7VKdExvea4wHH2ChVEgVmtRpJTzgG4+1e6DE0AYVXvnox7m+EvCdnp2
JUIZneRkRU2IH93ThvCuzt5GyRhxhkWsEby0WvD4jrybWYLf2Mi5enSxodVRUvmEWaApaXK1ObGL
3S235KUYh+ZQymXpywOADZ3qqZnfRflXk0IRxzkk+L0MYYJ0tGPew0LcgVL77CV6GKo36dDzJanr
S+7H/phpZM5U++IZqzrudPBu9yY8cWjiEgLgbq1TGmb0D30hCTdLSB66LkTdXfl6nttWikjkFa3c
/4d9vRNZMMVp4QOlJhNBhtN25E6g88chhcMQFpF0xZMuzXJhPldIaS1WcSnTJiT14v8pHVs+ZRCg
tL92MybA+9rEUa/SIPieDJWiwe0F8j/BN5YGPaIrAz16V94zOlrZuCpr5aKrOaNXh5AeaAEIqIt5
/vp98pM9n92WlBmGcWNzuWlEAJLpji4/dY3qvNLqeBmXHIyT2HMRHGvPUa0XI1AChryxJnQFDX8L
NrZ9j7B6FMTUjqfw40ckj4/2++PNzl5J+3gQT+IJIhKp1JJIJ9JJ2kXi2woXcKya/15BJjgewP6s
IIm8H0dN18ypkSWopcA93ah8O3OO0rBLFOwUaxhgUe7/GRnP6U54Jq+SDCcgCJHQOc16u1BTnqQ3
rCFDfk0FtMZWmpuZjsLRMUZIg4Ncclfn8uOKv3SxdCVEJNqk/P20oZWGlLmOa+TN96dzUuPgU1hg
6ipFgBJAaoThNmRjo5unom0b8lRLIJgHmXPvCh5LXRsUs5jetnWxwuqUGtI8mIm+gLgmm0C4YQy3
/27VnTdmrM8tnPmZB5qHmQ+KTCXTLm3jx+SIi/f8r9rn9YTaLXlBOEGa/kI9nFmuzHGKO5nwtFuX
5L8B7lwPCW9Ss36mvNfDQtLU926zoAwgNiYYhe3spoLy7ZNZvvFfCHqxGtEp2UWNObkWeVopnyfQ
tPms5OPL8yQx0ueP7FnfGJEKuHZ0SYI4mqUEEl7BKsjViUQ/mfNUnvI59RRU6Z5Co3Rp+2fPXYk4
zyEfoiH9LykgddnWtGeLPpRx2vBeVv32b7XCv3JjNx3p1B4tWLs8GeyDzG4VQSMh4+m1Ls2IPFd/
+au3nmcDLcPVWDAy8Yn1+JF7n8BH2k/k1y7Xv7QZ8X2/ZQ9MnaII082j2lFj12AjFxS34WRwMmgw
UTClPGog4XjPuIeBLAD4B4QfLC3ld5ObRU7kiooWHXhXuUm5K+3Ta3J2zeY47G5IEfh5+ePpyOMe
b+MeADlynxmqkhqUYG7B5F8Cz7JleTiGQHGuex4naRG1e63V7De1SV5pE/ICU7AKfNhZCuB0gs/R
2dATiMgCPfrgelkZh4oTznPmCLtzkeVNMay0u4i2lnl201fB/7RRREhmC8SZBVzdqn6b9Dy0unHN
Z5YsL2ORoxdZCh0G+EEoYsCX9IO6JXQiVQSngAh9XcCHnf7LtWkcFUq0yAsf0KwyqJ88wwthIfsh
vqdQxxACtfBISzkPVGca5Jv1lKaVXbGqke2nv5jISzVje0jnTtGLmDE8tvOvQI3uCUHxFPHp5c6b
4LZOP9HOcM/fDvlISkg8A5kkOMRpODV5F8tPt1Qbu1ZJP5IDU2VfLf71rzv8TAj6u7hZbkORO8B2
U6LZSTFtyze9PxzLHIZklMvzlGqVu2Ig0TeDGSSMVVZCPzO1Z3pZWYmFqfvdsZLKqy1uUX1wgZvu
E2YmEpMD3LFNvlQLOg1SSkdO+OsGoGdQKaSmM9NdC6unt96h8v+1eR7+wF28i2Z5YRhyTCpufbOj
eE/wwMAOGU2Qrpqti8IDNL+ofxEmRtCT77Rrgf7pP4hmxW3XgX9banmPTu1QD8X+Zm+iNwg4Zfbs
cxVYWHTSra0w/QibKm0ll4EYyjnE6hxAmQAd33Q8Y5pSIfZ9EYyuO5c2qaKl0JJr8RTc9OVPIfny
gtfggzTETF/oBMVQQuE1jf4wzQXVQBcfuk+K9UhfsdEVqZvX6pgiCmw7g0DilAkfV79p2qcMoTne
JAnHbOf9E6IV7M1XcTQc4SRsJMGPumAm5IUHLu/xZvhtRWB8cHQrlzn+zxVuFaQpdd3FOepCbVeR
8Mz7apKi6Im0TMNgCvYGQGr5hnKMV8ALWTMLrEpos1+tiTLn0DU5g6/nRK9lBZ3nfnsGHIEzhNp9
V6V0DXA59MfJuR9UuXV1elfgGjqDrHx9Tlt+iMYKo8xO5Ujuc0jDy6pZKv3RVIjGVPbUXgm7FpMm
Jg9F8tLKZrlwjPvYymeVYks4L6ClEa4enibKFtf+uS7Y0E2ylrJRwbLwqe6f+qnnlS0n2HJvarsq
GqNWjU52wPalgv5ZA1o3mv2jupf6GmZtRfa2am8T4GqkaQQs87Epvat5+39ZMrix3wBFpscLAGtd
L6CGcJ6pqVSyCFaLmyWWYNwnD+TdzFUeopd7NlMq5Vjka8fpDn4bjuAIQ1y6SOpMH0TmAbAXhdlG
pnXpO1U9k0jzboPfrkNAH6N1FRVSGQwQyxJRp1UCXzXPPITTTxT134tHypRPP/do5lWSoCx4SFA/
aI43huE4uKQEN+pbwJsy9dSC90GFRtR+MNsNECOvyT5BtJy2jRPAsOIAT6vxEktIKiwuLdNh5Q3H
OyOm5n3ItGLH8+arbu0DrzqCGLf4qZufMKWp+SbpmfjLHsB+Sul4A/kNmP9MQJdmqheu0dSUoG0l
lSmmCsjITvYKztvakWgYEzOPy7oTVdQFj+BPdO/tY08KpENrS2cKzwspl8ZxFmA0t+FydG0iiiDL
nL+qBf8aiFERCm0NBe9zkSrTd06IZupvP49k1U5lWvrt9C9mVgC/JFkeGSDJdAH3mtQfA6Yqv89u
LD646K2mLGYZ4i0vmIkVcOzV8xUhIxZJ6ajdxHuu8vvtSlP+4MlrLAz8jrchprbAGBraga/CD/xt
FV/Dl53adKwW7utjhyCTvG3CSbki7tygx4WicahL4NqOpHiMHIHIsAanwXYTsJPHN4gtjr14BCXv
Tey/WsuuNEsAj7tUO+Iy3PdCmu5SL4hdmSX4pWwRSZ76QwmN34KZZNLrdX7A31Zjs5x8kcBwGGPL
EjwbR9vJdPMB39GffDoDtg/qo4e9wsKnBrpfkaIPhZDcXUTEzsabe6Yw76+5DypAbBrdJ3RoPzf6
z7IetAtZVYC49a0169P7wuLbcrbKook+fBcKy/VxvLHFzOQbFXBxqdP5QseQf744cgsbQgJ0/dCT
qOQTsaE0To3KaZpJ7Y6hQtK+lh5MO7O3XNJRYzPyMiKFcJnMJthM/2etgl0uwroS4SigCnurDKjZ
wp1RzyYxSArHEvkM/cqpOSlv6GXkh70jCTJ2AUKDZYJxFrlxRSMBi4O599TWfVnvLSfp/OCFCK48
wiq3jbMG7Pc3V2Fr0aXjpEDZuAe2qT/ASwFsaWa/N2Ov0YYU6DelvwikZ0I8nFeR81aqYjzQ1ddx
aBLqPmUObl7nzc8KWmKti85cXtu3FsDMl5xzQax+z2mCJAq1TsyflwmvEFNGf1Wt6LChA2zBdjKc
6FlJKho7f6sjVkYiovPi7jV1tkNVKy8jXGGpMyltxBIFXCtg0FVd63Trh65cPz6AtkumrhGD/FrO
RnHf6WJ39xqcW2HA3bS8MxHZ1xxd77/rt9u7aHeTWkWWqXOE+CLc0hgUW3fWi901TgQfWp+sFFJr
kMLxrc8sTxlqUQHesDJnlcUlDbSvKya0B2lNbVdeXe5UAOjqHxDLUO/HfBIw2g3fFyEUiSX/AVo6
yh0TEMPcDHeUnaJALwwDPsLla4vCtr1zFGKtBzl+kI0S0FThuplMSDptuO2RvDE5inuxH8Bv+FFL
4aoGiONxARTemjleyl/5FUNN95rv5o3evzgYoaOV3KdrseuHRv6l+rHiRCfnoHXmJjGyg7MYBW4N
3j17ETOkswrMHt7Z/b4QjJZPVFmMrnSyOSShJatFEtohGgkMN1c3x9sdHqANjhKHHfQKu94rennl
IeKpaYD4V6fUz7fuAXjVRjMADdrCAFRoSOaJfzT8U4anIjZvnOtVoo1s6LB9dQR9OJum5i82snjV
zHGXV6OeHZBvVGJvqPGqkQNeJvMsxVEvuswADOhu0nJEo7PLGUlNfqffde600J/7i8TEXAM9W30y
t279J+lZKjmjSDiyDQXknNf/x4hmMsFrJ6tB5sJZSBkzlMs89LRomGL6JpJCxC2ZQZQgEgZLELtp
Eq6JTandPPL4Jf15f18VF0Qrr9uM1NDXpHPymByjBz9vyesmhDZAQmN+VfSBkT0q6lARWtZc1Mqr
T6NzE/h9Nj/hlmOz/RTHWspuqS4lVHZThgy5RbtAfklfuW6XR3dTnb2DXvebYMEj96b+9vGKaUN6
7IkKmhlwFCJwH7Kh65ZiUU7RnccTiGSb0cgFzvMHiY3Y266a0U5MxvaNNwb+99VLozUgM6gHGx2R
aJ3EWbawQy+x8Rf5p+zL1O9MnxpfT2Hp3fj+CA7yiHa06aJkQLlbWh7RJLTTKlsyjaKTzBW95cMU
0TPpSLCoQxCh7Bu5uFbQ8jadFF9q2kWueg5VvwZN2GixoAmA6OcxEFrrLKTwkP0OvM/W+wESZ5Yp
jNo8ox06kQPCYUd+0TFGyAT0m6BeXvXSn145j/uVqqSn5pj1wz7cW072sUau2bK8P/u4bd7B+mmF
1Hw1DP+ayCU8EHfAPWBthRbrly5HQpR93Xx1oYYtWDu0qG2DAKtYWxO5UMrTtN/LUUqzO/WNIzqV
DIMdXrViqcIKiHNtaea3wIYLjPPjpUMD8IeC+rThFuxo2zzZ0tU+xw8kThNTgTrWIW6gN1C0JQp2
TAaO4XuC2NOX8qE2Iji59glPlRyxyefvI5licO8UruUz1RgxBiCUgXgdla9rO7xx5dkFf2rOX4Xb
R5nO+gGpK6gXGARJCBHeHKidyAEDntUkpwGS57fCycKapAPZMAXLDGDAemCCoLabIKUnVHSyoE80
An3MGBZOa7a44LFMzZxyaALwKPyUwEW5z99WcB+sD8IMol0YREckmJjRUh50bfebGqC5gmM7lxW9
aC4dFAYj1MunxjgynVBskGR4JjWsg/QghW0nr5TiPIQtFRRrcc2JOIR5wZFpG6wJAug2yRZfWkSN
bqwR196cBo3LvmgBWOVdvQvdy7OAAAg1shYstQeNnsLaGcYIUhA6o15ROU5fhDeYvr2jCAVUIEwf
Ii7Z/t5G+HA+VHx4wcQJHBGe5F+Y9ivg5kYHJuB7RMb8bRVgAK+Ofv3QheT3Jvl/nH6RpOfOePpg
0fPFv3VQFZFx2+TxTPIz0U7Fsx35DDYkHkiJsaIHobUh5/mD29GtHqwzbxy35khKSJBX2Ufp/FHX
gNBNxzJwrh9XUDBpcC3BdpT7AWHakE6iU1D5CnXC2ibKFwNeouLadSW8HLV+cbF6ozuQp+3SXksQ
GVM0KMBu75PiEx942qcELk6DrCNgxq/TX9XJdBw772h2tf9XDqzFlwP+GbkEmnaKPf6db4LfqMzy
0fT9WgNXHrVUXz6nJCwa1A8vIjnMGEMnqHGc1DQ79dLxJrcz3DGJVZ285HSuklCJiMzF7qjkst23
Rz/L4pdOrbgPk/e8y2wTIIs2HGYToATJbZ0lAofQKxL5W0mO11waaE963rOTH0ldpwSwjI8TdyE9
DqHh+r4Db1VerUvGndkbuw3Qz4cNYQQ+94iNOWR66LlsDL95Q6Ib8aNcWfBYdMkgj9i9vJjt70MA
oEFGngZFG/uPZ0zk2rDq0YyjkHz5YYQPW09ISg73tNZDmtQKKpWY+XBttWU7vk80f1rMFFQC+5xz
VpxXbaJKrNA1eSgjAMbC8V6NkPUp5xQaedSiMPSzvUdKPOzq6oyxTvouftHwTw5aHe4V6QuYKpt2
lao6EOsENyohZNKV2cAAS+Txd75MfWreo4NsL0OH9ncCL+9tAHXuGfOGbpR/IRUGxF9S+KHqOfZK
NT+UDtEyfEcY2J0EwZIuowSQTX3UIGxydiLHWBUdgsabriXr6uKTX+UO9b7k9CXmiOx6P/R5MGqB
g+V1oArGzC18xkTzSOx/FLiAiS5jdIhOdzc8nq8pmiMtE2YbLJuGlOQDCHC+Dcc0OkQabFRTVkwM
9e3A2qA7+ogw7qpw/Qu4KZFbQ5N5QZlAlM6FrlKNPj8pfnpAU98C4jOWt9fl4pOAU2GHMY6rSOpx
AzJuWc02OC1lgRKBNZ7VMV2rImD0h6dFgKFzwGK62B/RDMThwoBkvyDJMDmD0GsDnwbmdFIKXKn7
yVQf2Oj3iGstX/Fu0cW9GCCDmga4Q6tGXVs/4CNL3UyckYkcPPD2j5NlEEgrSyV0g5QwIoVD2dbP
OojU1oO4o1DuMUCyrWmoIdWPyBl/MdJyHwOM0M+G3wvzNzWRDWG1GbZ4KlSyra7x68+eZQX2vmbv
UpJq0WsBA18lD7+644G+nXMEMAuWOyUbItDTdtD7p/sk7J/lRULC618PNZrzpVEQCiF8dIRgO3aG
irb6SzAPt+rXnSBmsWt/KOYjraOFAuT8r4ErfoDOmWY8P2DhnWKXnaiISVPdtpu2XeRmRDxCGsW6
WcQOI6Osen7K9vl5SbMqA3MQKGwHFr2BzCyCaljBP0G/XUXusWCMKGANifszLLzBS5LI0lFx2dUm
BKmcXhVxgkEZNCjnYCs5rhwgb6hA9tcgs5dnMnbMGuy1zuFPnFz9zp0kR/ACyFBv+mlRWbEr7dvO
ywKpgpUS9y0lssvaj0vMhir802V1WuVaRAEYs70IRwJd5zFcl7g6r8wwHtfyX+LepnjrhnLI4VRM
mvNDDbGEnGNF6z413E/Fk2jyU3YpmAmJ+sRuqKNyWuAWdeLE7bWQg2u+a0SAEAiqdWDvYq/VdV4K
EstqfG2pwwDXwsYdnMHvc916FGY6GD1A0m4ywAvnWh/IX51zX2f8uF0kj05qcwtfc2Pp6/6XgT3m
i3gs+zfH5Z6CNFqtuK7+7GAQ7vfxCuYGYcclQezYTca1dqPQEBVHDzA9WFGr5oFpO1ztyGgxc7xB
K03Lp6tvTSTF5c04lpiDtWy90xqgt+dRwESkzXqgGsgBEyOp5UeNhkg1cSql6lJ0L24c3N+cfrjj
SfSomwQuGyZX7IUUMyBW3SuOYEzV+Ab5BK1RFZKetvryw/eXuJ9L1/uR6aH8Yvpgv4fApMKms8ES
8i+XURtCZvPTxE8jMMln5f3suxvb9cDUPNPsvRQQv1dtLCqNyq42G2DfHBh9IRehXpc4+CClA5Br
HJZmBaQA99ylc9+69cV4CXmbGbrFHMZLdFtMFZ9Z1ivfC2HDIY2amO7JKAMGU6wYpptxOQYRryik
oYpFSll+thKmp+++UPtJZqcMl7lRe1AFATgi7VQY74ZpLfPiwnsZxMaD2F5Gco+Q+XMeKdkSYCi1
lQ1gvVatsx8b8DVKkGYHOlPGV6salpMQN663fqcrAZiXdTzeU6YOOuxENIpWexwtIsoj05AboLFo
mc9GFVv5+SSrEaptImYsqonbrcsRHabvD3a1IgXzExTzWBUUbc75XAZBAaDTL2Dj0bM2m+KNoWpm
Np+DlGrFvJx9uPajgwDJSjhjKsGskVtBeawo1NULHSCY+ZPLwFNv5cHoGv1cmaB60rBghBSbA8b1
0fGmjgigpj/1BVXc8JRQf2l6LCyduFeHvZ4eo0VQDbLr/XKwTw04oPwbcAvgIBx3PjLLHmTlWX8k
4chU6DzOZ0XZq5e9w9rztWoBAuncEXv87nPCHDJ68gkqVrc7jqgeUUUQ8PG8ezhozdRurnz7mSkr
RG6b4T/DBTnJXF3Fn8CvNHXv01oI9pnyy7VMeFgAtm/xCWL2nRLtzMSAxwyw84m+x+v8YNGhZ0LM
iYRa6iFhAMRVMJJ+ZBuuurZQ2SOrw7eFzGLhqIC8H5MKvtpRq2KgjjNrNBBfF5vNIIjULVbgoTaa
PFvR51FAlUu1UClOyiZ+DdKdfB4U11IcDU43z12Zyx16j66jEZMXMcOb3xoqZc4s5hpTzfM8dGJ2
5prbiCebPALj7DQYfbBR125bQLppzMiFCqKMCzSvh6BD0V7dFAWI56t4kpO6kNwqbmSpgWrft+8s
O0gEu2JWbiThavEO24bvDfT+Zr3Y7xcCu2MMQJxUFVobXqR1Y9/+Egc/5r3h4nfMjeYfZjiBVLdU
2gftINGscBxva6DPkGK5W5/pmSNX7lbOgf0UYQjaIAtqkjBrKpdzvDa2DXOp3Txnfy8fFa88QpP0
cdjQFK9fvb+v6ypV56SnML5EHlizLLPxB1NdRvwvajLA3vhAZqQc6PUtwHh5epOD5IrGzVwpWxVz
E9ubuScHWStjkVz9TNSajCgWIEA8HyqOt/uf9nnzjN2VxYOmh8zAbOVYMOHHGMbaxMqZrYGdQXgz
/f92kXlvf1RVzrhVjfXzQ33YiBWNEzqS4DlZebJ5iAqaLGbeI1kS+D+sux6wUQVVn+32IMkaK1T/
5NNfo/8EB97Wr6qTCBChIEXEqjOlud3EIHdC9nIdHaVrZiKoeVl10yYaFR0XEh76SVgES18lZAq4
hSTGP04pUN29ZlujaB0BGrK1v6lTtCXTV3ueldfJR6kU/wzeIK/DhTnzp2DaskHaTu1dg69ryiqB
AVGinqN1Ic2FZzcLT1hcOb4zYh5G+MZQgweJoBYNvZtHQ2odJg77RS6PvCbEDu9edBdVkohjhyG6
qT+We7AexgGrx+aw1OIBREnmUeLQP4XVHL7CFL0fjjCoTU52gXfocugbtfDUQYASf/EdfF1HHscv
D/WtzyoqCTmDXEMtHKePrTnIxnBePV1DCfFAK9K1iYFHyUer5kU8cUC1nmfGDA+kvsjEEzsgAjok
OoGuqiN9QivkMD44yc/ZDOYGlP/toOFb8/yTWqUxd4HdqTz7T9Wphz2Qe/2kpVpR2hIXKxLRCbK5
iQIMChabd1swI8uCfJqZBGXQdgMirwrxDhIdq0Ampm2XJ6XgqpwfBEcAfkQnhw5mXkSv9Xru0jWb
igMzGeftkmgP1HMglo+37LXF95RxSMQcPbaGhNJbqmv4C8k7s/bVuRrDjUBviymU4X9tsjdXRGKc
FGbA++TdbCmX/i8l97fQmE2Dv85zQlG2l6mbbX6HeBq2kEAB5PlWUBx/Qa72xEW3gIscA8LZahZj
CEVAHe9fALtuWmvXCpeA4WHDnB9ehIKuZCaAK6kY5VnpXI79UPmsAQWHFiWymSrbsCyYBWmSnlbB
FPE7CX2ce5Kj9XnuHKghQZPhiF0ne8e+VXVcf+ZXNLpZ2AC4/xDWE3fBZXBO+Cg8N77TRJpBsFaH
LhF+AHYmHyRaCBRWQAReU5i4xNyp4wpxXKZhtCWMSr8wmGkoidw+EK00dRa5HICj1J2NF8C6wdFi
YzNVtbgyWhFWugVusg1g7fGASkKVQ768c0G1GvFm0ZPPIuhXfnd7DUpkdGmTFBrFL3d07FZWBWsp
WksBipKSvH9vAys3fnmHiHM600TkqFBSvts+p2IWS56u6fxWcQ99UotbSH8QPHL8Zx/wjDaCHFD8
9CtUWiPOsyNHpBtigImTaO2HgNSmgiNe6ASY/XhMHwvYIZpw9o0YHAyEYspnno9q9ZQ+jJOQ0oFb
EAmXE9apAYNKo37gxe2sihayt+6XKpYghgnuaMZLft+Z7KMdJ+jbzI/DsKKYfvDju9Vph/XssntM
vcgUwYLBJtUsyOvVcXAxFOE9BBkawWsiBfh/C8jTdl/5gqn+UkAaUUZezUCXbr3Zakm4dePIJ8ik
GRPVOVTV0hm74wIMnnQSLvahb9HnHQsnlx0dHhpAFdVa7LCh2T1anuJ4bv/rcatFu5SAD6//ZKOp
651lOqI3dTCxKt6QS/Yx6nrLIsKRPVyLz95jqtmQ/ZUJjChqUl6fa1XJamnQDBOu+vW1gyie0c1S
o6g2URM+u6jMITwzdEgHFfYg0WCtbrIG+4q4P7dni+qX5wH63RAdZusOfzx2e5EPDeOsveH81P+e
zacAmVN85zFV0LUMer0kFyAyBjXjyuaYtIwKd8K5csxSMOOIKGZlJXRj6IwDZ4KPVC1QWhrAiRD4
00ZGBC13TCD4XMbjl9wf4hUyNzoyNl/TplcjM8C7iTrBsYq788v1+aXU/Qpx9qToACk6h6KbGfdt
9gQOLxVHZKIJXCssNoyzWuOtA0YeS/n5cO9f9AS8OjC3HDRmbhsPaysvoNGeu+956WVVIbknB41/
oMCCrFRQShnEhKwdJXdQ4h6QgOGC7lQB8rkt1oJpLFqdxN/ZVPYG7HsBbWkDSHcPFoNPVEBJuFPY
AGtfsyDjHFPbfsVXxJyDgbT9ZLB89bZfw0TmO2BTBMz1nBOBf9w0wcdRdinAYGCwCqpyQf1/dTQs
iVGyh6nZpMrYeuIXOXmQVXxqc1wb+SQIrxMYI3mEwq+clEgpPDHcYREkindXsye4vIbxieMy60Vs
4f03U10qjmCAM6+vZnhcbt3+CPwMQNKvJCY4D0STCX7MqTl2qgKJhXqKsCC+Ut+BIlL71PzElAXZ
9M9EiGlPuFRv+X9P2Sz4g8pLbb6F9BM4niJ4gfKx3CrtOIS9BDzYqu+/8WKASXSJ4H7EHfLmLJn+
SDyiu1utkUc1sfDhKRcrerKwL99ZK0Rx1Vybf9/xQK6bvGzbgWjaNspSVzlE8PQsuK7KT2JylgEO
YSsCZQDUAIhxPzYNcZOzKsfQz7/pdTtcmQIvB25jIcKZMRFWEM1B4Rbz9LFwpJlgn/bhBSPGv/mP
CGQ/PFFiu9cBk/1ShHnDxawdFPYKohfbqvgZj3CvSNA32EMHErIBUPB/6Xmj2XN2ceN1vl+40w7Q
CVIVrC+VkRFV2lb5YNEuIZe+sWTZ2KbJK38nOk5Kv6L6nd0sO0dhQ4VmQStx2PZERCiEHXe1UkUw
nSDFHOQXOoR836kp+24BHAAYpmqHSxQZiJKi/DTofj+4u1eiuQyFfOLPQ0kmiE0cR9/otiyUoNF9
RXJ9TlocLnsKkcE5/DU1VzAiC2GwT7o8hs+Zd+b+XEHfgSHNa5oUkDKD8NMoVAwv/MxBFQULQ4/G
1fRvUJ4Bc2OP0tuC0t1SMq2/XA+FSucNfUigfppsKo7ZmE/JVqfqlrXw5JWwKqnPFWv2nx11UJvw
TEMPebaXcXY6EJmuXIPmFC+opEw5IrM4yhJdjSg846rj74K/m9sczkchsy19leyej802ZjTGl0rd
y0texXY4luv1bgbVDiZ7yF5mmpi8riTTA7GYAhXJ2A6mgCzjANgVp3XjxyeVNnK1kffHBNHeET6/
XUV1OnjhrgQyz97rP1ovVHeeFNqKiIWJJk3K8mmO5zU3/ok1hE7cMYW5eidDK+piYRSUdF+SHHe6
sPCcAy9dopJTJuU1V9wmU6MilQxL77u970GZQDFmufMxZNhdTUPH0w86TvkhVitR3pKiBWbVtJRr
ykHIhhOkeRmxywgYOMBz7VFsNoJQZx1i8PzmtkjoyMDDctvHpQZAMVgiVYhLuRTJQ9py064NNQvp
nkshXG5PJCg9PhoSJpEt+4oTSk5HSNlr914VgeYwonW3e6Os+SzLG3SnAwhZcCFp2xIJIKB94Rhq
f1WgeNPfQyn7sTmsAZ2HlaXtMAHEqa6hp7uOuCJPkGb6UR0Zrr6xZ/8K3OjQx30SrNyfho+jVJlp
+EF1tCuBVcV6LQ7NxKjEnJ9HFtVoPUwm71PlR6SF4/8YbigCjgUo2c3j6cHLg6mcjS2RExUjPa09
WVku1VH4Dq/PTOZzRcfPjYSOBmyuutbMfJlRuosMntGJiWgJxoVr1k3DjndkZkqgU7rAELnXf47T
zJE1NngcEBWDP6bCi0mfzaLWhbidzp7qQM0OsDUj9EDf8J8w2AoPZLt8xvMoKnz2qLEpzAgyTUIP
3fJaF2bKIvHlu08edN1wWHbuvlTxJMkIti5225htqwyZ1d2t1y/LVlOmFXr6Q1JKWB6nrUgKTKqG
sKVzXKpTQeDvxNff49Ul89zz7geePTknUgnqgYfPlFEaKd8iFYt0tKHx34UXsN4a2CXsd5iKhTjQ
Ml+b26zuzVkq4WaGcRw+CvazS7FrjgQINb1Y8UEaZe33GGici4tLMmKDkMtXJGbgIUt8a3wBU1DB
Bjj8DKObmeZPv9lYdWjgQDuDE9wx8S9Lnql71J4hTsxwc1E1YBwyM1cuud8+jVTLTQp0D+VXKQw3
ehXLGpy/gE1aVj/Rmd/47U76K+xjPbnagDAtbzZx4R/eJNEw8xImO0Hj1fOKCD1lGPmmZ4JSwuGY
a6/vIviqJ3rDXqud3OO5nLYFNILb4YGnkkizy/y8fafoE553ZNwdSCravs6L2BP9Z9YJVR0xS4Ak
cun+0knoxAifaEB/PH79ZYJy2Y///Fx+QTaISx7JbGp0sMEDzWeZ/GO7n2WIO8r5rf9bVQj8HpX8
VJFnR6cm3Aqn9vw7etbrM2DB6yaSu3O9WC2aOl5go+aGXAzUOgVF1R50061Me+Z0B0oNcAyS9LRf
sXJ2UN+PTh6HhKF0FWV/VmT4aXtyey03E4TYWYN8jsK2xqkPNPZz5xD/Jz6JAPrMFD+4k4kFmFlb
QTihNU7qr6XcbKAv07JbwW/TerUjVXK5uI9ItoUQc3rSNnBIqXOJQ9c+K3wS0faIswqTvDOmkoxE
d7tWmXR/NLyV0U4WvmX8h1lr7yuLCIi4k097iWk34cyOr8Ur0cwv07hJ4F2vEK5HGzi6hYSCWRjE
XJV1TQB3sclI4XLSczTRvFfQ4rMaZsl26Gb/e6Q1od9tCHYFfhtCJOt+j4BPK6GuI02TuU3F/x8H
lCpdH7hsz2j5J0G7F7jMVgFUqlwf4z2kcSfOC4zZK9kqNheFEWDbDBPlMFbheQ9DERIcTpJkTaIH
940tu5rAq71/1RokCPc/ZTA6369X1ISDAtwtptRX5lBDIKRWmT6QfgoWMD361yEW74pI2qb+jnXN
eHIRLecSp/sWRVfg7tTaeAwxtRg7UZkdoF3LIyY3Iza4s7xlGfebYBC1sBrWVVHzjT9s1sVMguc7
3SD06KQXQvpY/f4djVlUV3WyGQGT1NH0CiA0DfEG99DDS9jpLTSOQuOFRDu14DBs0qQc3UrGku1a
D6Mp38ZOYelUkLr2Nhtl68QShQbeTpZOsR3A8VTnvcPYQe7ztNNb0eMoln8T5JnXv7YG93zcLAbq
98SA+NkM18si6lG7MB8mi4bhGPXiUrjOSTnwTay0s7UoUi85S1ZTOie7LQCMtlPowo0MFipbr8QR
muDQnWGRrmMt6VLxdmPw32+KshIemjd7uF+MHlpy6D1bGM7I+XX+d9N3OZZEQxRYUvhpL3hyFWkk
iW7+d9IhXnWcVPTqWpXgTuwWX6SSWfdk3W3DwFvDaZHNLKFlhYFRPwGlD1pBYAfvJUhdDBN8/MXo
0ZDYDCKyvBm9Ry6H/qOYq8tiU/92k5ba78MIzO+NMywwjAi9ynb8Z60QhREzbjsCRHMoyiCGWrRB
FOGBh3G3QtlItaaTn1YVB8Jg9xqNzHFnnmgbo8E4dyL9fa6cEaIWO8Y/++4DyqSzlLyrsr0IIGC2
1FCqbjnSN/DuwvWi1dtGCDxDZJBSGjL0PTNUDfsg/XLgjmz0h6W/q9zZvV8cMj6iVYb6Jj7GEo2P
5ShRCtfXpwAiZYs6QRuqNb+cnsGmGmW+kNThcAKzAaURLl5zUefZIqnShZNFIqV1kuDYuji9ARRe
h7KhnWOZ0B525x31eN4cpS49rnk0/gv/b5/Dk3SQkU5vMYsRgbrjORTC0AaZtwYWb7m90TZENNOh
uIlROpK2KZ8VcmXMbwf+jWj/96U7KfdMwTWGgZ3Q2oe65FjJRMrte6yDIfWFcCkwc1CSs7/e7+FY
HAmyl1CiBCOjC96sBCyHnGj/IQgJn4tl24mx22rNG5XDOIGvOGJ6Vkdb7JMPua+S6g44+NfHDflp
TLzsISyWv5bgExxah2SDuIZ4tBzBB/finHw7ZyeklvL1DSTNNrhFcARaJiLcsY0t/mxYdul4VgOv
V98XZBl18/Z9O8sA3zfALUV3I+ksxT1FezXLLQEcEgXXiKDFJ6dAW8E0mlTrlepiO9bttPfFPlMR
AsnautNCG/LEGv2q7zv/MCRcZbldbqrlLLwCXclyXGWFkMnfO+mhbi5V36nOltjAjyIZ4U011hPU
IWgtU1lvRO1jzTzIzKJnaqBmwt17//VNY8ANdPSODDRTfhHVWnWaBiEO1vq5I54DboY2tt6MbCwo
2uOQ/vQZhMxqFzY9zo79m4b18Jz4LDMV6fGEMEuijOVe85Y7K+7PTY4PXGbbAWjQhHVpLPaG6ZDy
Zg61bRM0kWJ+bJOjp7JBeGN88oYyDOBB7pyqHUDG/Ofbkk7dmSb/4IHGMXcj9UEq2Hdl80tM5ym9
uabLjdWhvwxXjKyQr9zUA8s+Ln8f0SDko2DfBdH++SbuYOTERYL7rkbSreeEvn1RZ9r9KkbX66Gb
rsVyWbg9/etJT35GyY0NUTu61WFykWOgdaM2ltOp8LsWoqa4QsYpJVLfIKhFSB1jcQ2fOPzJhdvN
HA8o6cKfgHpCPPOhO9DlpCanI6VnakY9gFo7kO8eP4iirwDirZ4jWXfOBnzD/6gmBDTa5Sk4juIV
SAnwC5wWLHYzIpcQkCWUeIPs4/cjqwAYNf5/ur5G6N2NSyj5uK5d9NLRz4anRxaDOri80H7KmPXU
1i1sG+xlAeYI+gO5gpM6lLiZ3bGgSjmZ8+skGs3iF3AwZpPtkMcXJEzYt0qxnaLWnTWn7y9TTple
32M+85u7Cfff3A+U4B+LH/wBiJMbCFOw9BchtKQQwviywUSJsQQ+0+pO0VJTsFxSJN2ZE9TTTKmb
WwHmRDy530UFqGLx4zTnObuutNL+fEmCrFU7fWf74c74khxQyO18p8jgcOfVI/RwayP1O/Ming3f
efkoPEJMPmyp6gCwnDuohjf5tlS8ROdOjEDoKGJtuw+Yo60z4+gIyz07C5hWV9PE04OeiH12zUCy
UhOeSnQH0HCbiHysT33BEzi+T/8Q4k93BnEQ96XMJapxTk8WdXrFnOn9ijGOFgcpsmLPW5C35PjF
SWVjqQySPdvMVAj7timfeThIlqMWvzWnqgZRUtpMmP7IZHQ70fsilSmalb/lNYFylhKgHD9ceJbj
1nKwuxshBBfi+UovxQby+MJfh3mnYSlQmXnboG0iejODncC888RFoVuPuAwQgOiHwHnbCgt9NWrz
A0XSxxkNMed/OaV3suimoiw6wsm/Ei2c22L8EDp5G0mEXWuYf+SWEC8bCagoodkRpMx8XPm5Gq7D
+W2hOOH+BRpmLMNxZkZpaFrr5wYZoaAQCsYmsaWS73pIEq5HEAA2kTjAq0NjtIJASoy4vwYOBffI
7el32Ke+Umwti3Vwndepbq88IA48pTMvzS++3eacM15qBGxHLST6/Ho2r7xQ7SnKQLaQQNLnel5d
/lE+MdDL3Nc4KmjUv++14ndUfagTXLqeWZp8Tl1nx1zaFXxsvOZZ4qNVMwuDBEw4BjraTSVxEMYh
veTLhmbIrOOR3m/F//wHlkX3adKq9ZWsesNLglkrbmcUu3H6OM0BdhxiNUWSKDA5AKEcMW23nhXv
/dkKsxa24plfLT5aYnvkKGMvSLRp+uvBh/P7OfCdnqJiQ1j6JMHRxXwm4XH8msxBFg6FlUopBQ9I
vYGWCSmLS44jH0cY/xoTYVaQ+a+oQLcOOOiug/JyEB7kRbGlq7hbltGuKv5b5qjbhsiZR0qQoT76
JfGMBNmXLNgLurpONelv/vTT6onrlejBzknJuggPtZX16OHKyawCokqqUSsQ3JiKdd83QJtlduSx
1erm1A5qk4CTGjSLFNXa2RC4pxyilwMlZog0mniF670BnlKirZ8rqtgx1Ht/5DU6U7U1WxwhhIR7
jDzZvl8GC9RI6tY0toR6FrY0Tst99b3xA9JQYQepbU2TymSdkDfwPYm/t0MgkLqvn+hXEgCi8VEt
0M+aQEC+2Egnhbxb0KiuHsu9vDFOneaIDgYfKU5yec8Ix5EYkN6pfLoU7Qla0AdiSFsUwKp0qKXR
MlpUWHiv2ZKlRdVH5tvA6nsE3a/hpI+zQPRAoYwntzpmUMX64pwrV1BKi2Ed8znAwcS3fCS6O3BD
KyJP5ZU/2o1bd0Gp0PwRvpSlMbmMwnV0elQS238LGuDh/S+iTR5E3KOQ72Xw6lKExPIqYUv+bAB0
HmVulBan7EWjkiYCYiUa1+9kIBobn7AQxhSB5jycy9wi7hiFWeKJjdkxuQ5Y7W5Mcl1E7d5cuH2Q
X8Q8f2XQoycYaLP2IB8aw7gSCY/R/8oIWBA3Ifm9CXTcaRnhDgjLSqr2u93/LVRc32M0APzuK1Vr
dNHuOC8y6RjdBBHeLYs51XKYB6ZF4YEwJZLNSxE5AO3UWb0g23eAHaxe2LhXezLdIC8UjpwkB2Gc
xBHk+BQgQKB8QDgI7OqZYGbSDszC6Sd2m6ywBu4HxzRrXIwhHoGWRV6MhfXPwT6b/tfxT69cJX3z
FuytPBvvBezXbcTks1bbNheJx6xksh+YLnC9HiXi7H5wSYfYmXRHFtyVue+Xdb/E4NieRpkzMR64
zTBoRz3tGy7rG9Od4CUNpm88rZe+LXMGghMg8ZpaD0qRwlgvj4fXzLcmpPt2D16qSZ6x/ZaZYAuv
70W5uRYomLOI2Cjy4ZBRrHcr/8unjKSZcVo67GA944RvDVzmgh/kp5VtSZxay2r9Cv40spvSdoA4
I09ewy5g7FT78NMtDwZvD8KT025w/M0lrXHTtsO/etj0qVSZdCVeTqBPrU8KAjBfXjnRTu7Vhu43
uHWs5UAoAwDwl+wFiPmSRhlM08RW36N8bSexjFFUr1WEY85o5+6DCxamq/uF7eJ/jSJ9RaZvEgFP
Ejr+J4i1b/F6IAIm3DKGXKNPqpLbS49Wj07E06advXvtTT7nwYxlIfb8kI0+NH3UryMKRDplKBY6
gtuW7e05Qox1dKm1gt5yXy1sdHC09S4diL7qc1cKxN7u1xd8g1JnvWeGfrNPQ1OH8bFZoJt2icLN
UwbN01lktvPr2wsdu+ypu1ABGGikJ4Th5MmDQeaxXxtyI8IQZs/biIB+ZRSD90XDGMbJ0PXTjhzD
DOFjl9mietiJxwZxSaL7G0nPrHfC+kq9dUuf4g7DUd75cNH+6G1XmJqbWDd1cI0IXrgl67k5OJK2
NKFaWTk79nBzoDHkuOUdkD84f42wI9u109eZOkvU09Mmjf3oQq+OhQg2wMvflrSN7/Kxjbw01bog
4NaaMflNpcUfyJVgU37iFZLOPNPlsrXXAX3jrk0IvPIfohzWvxCUU78yzeD89ChHq8u50bXperEL
mkdPsefIPOOyybBV6qhpe/fZmlE4nN7uUSfdSM2PeEDfFy8eRosk6N1o6VOKoi2eBwZO3zcG4GQP
fUy2VeIfhR0BLicaLdNhE7ZmZoRNiml4f/9rw/QBAI9nzXO3COHt0PRd+Yi1oHh0t0MSaSMmvEDw
pTnmPHThsn6jwl/41YKwzhLXeFXqcfKXfUk6LamiqE+uiqPsG/CLbriXri2gUApNxMJqzPOfMxE0
IdXMcF8KXc/5IGw5ONKwehIzGpLgiiQTMe+4XNK5HV54Tf5up+6tVhrav4tzVo737LV0R1KN2LbA
pOVwWc7iP3G8rousVZywujTv4Vi3owWWf8hDaxj763F/57Dw6uyIzcyOW0+rDkExbQtlmFI9dRP2
hwQwl8Ia+0Il4xNEQVsI9KGI+MQhtVuvzkqObrWBJokOXJmNRhRwjK3YhFlqu25XLOoMduHWlWUM
TCW7cS0e4mudQSpLs/GsFAbKPBfBLGzIItsDZvDJC75V08UU4d4MwogCWGvjLkjv8UsEVHMR4RQP
LS567Ux+5s9eFiX90/ANAJhtj+1Y9l/9B7+LGGJT+KmvyFUT2ZQGk+UMdsfa38IYZPXbqR2CR0vH
krMFhev+Qs66gu+rkuA8ymFrb8phJ2LfubRJj4dmcQCo2wHK3xID9l1DhYNaBkBuR1Hbz2LI82c9
a+tqahcf4HIR7KAgb4w2WFJ/6Iqi8jhuJBjZqLOeDr5GtAQQFo5On6vpmN1GPsSdVJdTu0Nge+/o
Ze/zpG7BOF78EUfrzNACiS1cx8Ocsjy8E8/UKcPEA6c9C52ohcvF6UcGC2XOlZWdw+n4Lr8RMzF7
Vtglm9nctNeygGqf9WizJBm5++IMfPh0WHxj/r87GQLkfJIYqu8uGyyD5g3AetIlJSOylcBdyVNH
C4XWJmE8J85r9YZEtAMMgYv2Dt2XRWYOcLVwX5zgNwlIrKYdSYo9qj9aB4jr14pqn3ewhwNYiw7c
Qr1ev5JVuPQ4AX61JKTqTNRa/gfte8XZMC7syg/73nmXBh/NFNZrPmSSsMBGJthhH1//vpH8PHBZ
P222NnQOv3ftTUDMyePyiz0bdCdZ810p5n8cj9Id2I1u7q57KPowfILDd0/w6eeeaN4kEnpZWJS+
CwZTHqMqr55uOIO0bKd1a8NP7ObX8Lr2PWffwwPhTJgrNkaVYTuaIh9EiqEVsNRdOr9+vChJGQqT
hC18yd5czT151nHSYJx+OiplAWFOBO2W8V2fGHHqPh0FxRm5wNay0NuYG300waI1GsA0hcWfqNDR
9DsJbku2nF/+Z9P6If6/+53rfxUEq6D593q5TcKUziwfW2fiQ03wjnLj4LcRFTjbt48k7zrlTfML
bxlM+34qJnkOYkdajXqBc81xqbYwdu9zl0Hrh1/tZDIld97TnvBEcr+CltLhXf9xle7sLu2HWZUw
0A+8sSkGouD2EQrEdX4gBlS7x4HUB16j5n7dF5KThJF7jssEmLMyinqjffJr7cgotcFDVyjLf541
RkY0/ujM0WsiP436HKwFdVYnM52r54D0/E0lGPxpmCDDpfJ7yuOnFHbHSDngo+SUuxV2XXvHax0m
ewiXUVzaI0360IzKZvdx9nQiIImlQJYpW2pobFQjSHozAw9TT+WftDiyLKwAfitGzSO5QZXKA/4C
VTJlCEx6pUdrijs+BBdbIEBHorMDFLo9HQVJhVAFjOrKzUBdKQ25wifxgWSMGUsjgiZUjZIDTfKO
iLtnrNsai/OQmBK0BoE+l1es1r/H3KZkMoa8GA1Ck0y2DxKN9b9QSx8XXOUMYFVoNTh2ClummiXh
oK7C4IBe98cz3C4LR+tiA6LrIh2dWulDRFBqfTPSF9nDX6Uewi9Ve4eqUHh+CQ/sdJtelXIU0Iwn
hEVyjC4iiIlnUboKD/VI1HiuFUKh5f/DvLnl+43mkp+6pnaopfRSRJgsSf3lN6hPoL7oGg05NL16
IcaX/eNqe3Q5niNwGTweu/j6WqCR60si8gxewknzGdLrzwnJ3+AeTRI8AXQozSGadgbvZpQGp5+p
kxcSrcXcr6xr8QXUoXb0IftP0Vbz5k2rUGLXtWv+gyuJ9yFkp6kBl6fwAHofVGYy3lWzQcxrFxfz
L0kpDPZD5sB+wzV+OQVc5AKW4CpGtAYbiCxrh2muQdiwFc69+T3lWjF/aFIfYbocdL6cTT20wTUZ
0+z6+iENOLc2KhTWCdP9nJ747PR2CEE64oDfjMkQFb8slJCgCvMZmK0+tUUXbSaEj0j/awWPdo6I
xr/lTN9bJXhyUb8sVNiTq60/y/L9e/M6n6m8Q3bkopVro+U3RLla945a7ryaJAAWSiZF0OdGEGtl
X3HwtsxRhTuSP55PivYe5zVAJXgPk7cSbgTsz0B7+UicLbchi4DCx2rAzkcCc79pL319/clsDU/B
DFErE+qs71HC2nTUN10Wu9U/Y012nKUXYfzxUefl0tVOza4AeJURdZoz4xEsmlpm9Y4a2pk5EPf8
WPQpfwQOl1WRZffwfEdEcD3u5IPc0YJJk8FBXs5BCPGKVvuj20RmnZpDNjTUJKnUGvTj5tiQBWER
Vaxgptil00/+akwoqByZJvTUSG5h1NTdbSG3pHlucXtMLECkx/KrO/Ovqfdtq0OqYj7RITgSGwuV
XXi4UlVxuH6Q3gOZXpNMCOgos+d8Uodgjwh0sjBHN02LD7WWGubx522k+du1zwveIdqCOBEtFyHH
96PlknRMZIAoz/x4qliut9/A5+jXrXfkSF4pi6auTLX0Wj0yTd4/G5J6jk9hObtU5g52+kJXq04p
ncM/MsXWj8jfO/L165fGkgmSuvqoBXix8lD4brFaJKJpXGJwHoQdbrKWv7dH8vRzq4ejnt7L3sTy
LPupRjNLnVmMXgBipcR2IVHGajvXb6rh71YV6kme8RMG0i+ZtfQBxFTv1cgxs34UE3nhYXWUFCKD
CLnFwKwJgeMo48IMbXE1TLiW293ek1oG9nNbg7/vo3ClcgycaPwCd5wPUiMXRfBHqHcOZKHtRa1Q
8t9lO3lFuVyUCthVbLC4MJarMMOfbNnJud3vJNS3bX0dBCkJF497F8jEViMd25RUFZN5tb+syd4C
fkyRQmEq6q1LWYCKen9zr8BTd09ciEekuZISpyx7OL0+ct10aIRjaJj0kY0jP83xpyL0flTt9tY8
h/t8hVNy/RhXNChY7prOhUROnJSZ4AWO9xofQQZ36D/vgfORtNfIJ7Bp6WoYXS9rUkDdEa3/Hdk9
y+mNInZW/pDIP/vHaD4P28lgn8Z/4mCgPC5ZEkItKjc1u/pS+uTPLzUKjyKHPQkUmWbJuP3skbWu
F76Y5bKem9YkU469DojmeE/lIwpTNUjE5di5T1vzMK8y2sdkLLBpPeKoOkqvs/6r48TJuDXd3qrB
oauZpwmtAWSqvkh8An79d1KdSKbBsQuFoieN7GjJRYzosShL7/GzTZ+awAmdOrBvV3Q2L1bKoUj5
mWp3KAsjAOdJeH6n9CuQt8SE0WiIHgmVF+zCLZkOvgcPF1aRWAk6HCGaJupnjhKpBQlm5TCDoIOW
AStTJV5JQ1xSPCiKMUV9HrQeFqBg07ch/3WPANyVL1ThJGOkbFgml93AYLxEV8KbvVB9RCUqdDXD
zvVcHq4B//DV+SpmA5dQk/v7BLtFZO0HIHWhq8cT2RhByvJN8b823fkoB1W2/37ge7E3oc5I7i7T
62XRgo7rbGD2SrR/8jkCbzusolE+yxO/oEXkLx48hD9bzRnb39K8CPx3kUxQtys5jNR/VAGAbIcl
hU+JdE5cpKkpVFjQZVfOAwkOO3cnX3BPb3nf7I9lJy0p8u0h8W1dJvo6YlBxqlp1ZeKgxu+AhgE2
td1nI6ejOGPoystfsE4obKPaSlS/j6WMoi9GNmh0m+8gcFpRyUhSsSPJ5MEFsNsVRyxXDXRJ7qjk
bmAfqI38bKkkyyJvKTHB1aZSN45OJkWZNjFi4AI2a2fd5efPwNAorToqXLwRKYueU+wk07T/5J51
TBkrpXAqx20eXyPqm24grI9iexPN8bMbZrusA4zlS+IMIGjKStz1MHrtqsWfrmsNrjTu/LPsxlAk
ly9iXLtlMHYv6qVM8buBW65cvV6uGVMU9/Rdyd41BkM0C3u3DXF5PAh+JqmC+j+3db/4PW7fBIL9
ieVZ/k6CDCVwJUg+PjNNVyS7iwyyYRotKFCGxnwOae6+OkOagXXwpz/4HMI9wEYsKkBk0Gv5Il+H
3Nl0YM8IUZmArfCkOyoI4GDhBFTU0j22sc/2d99xLcYdAh1lMN7zqBbl90qmuNBRaLsfnf9XFr1h
pm6mb+VVtdpvRBWJ30bLnw1pVkMD6+Z4YK4uYtNtCtK+y8t17iZKmO+BYahHPLh61PTeRTZEHNGD
oes5FCnu02FXsRRevxnFnlcBkoWoGkrWKth/HvPWdLKtviXtBZEPaO/l3rgmE56MhB3ztsvsXFZ+
lUxxXBv6jGWKjP8MxjvclWXCcJ72Hk14CGaSz9bvagZtvGGWcmZSvCAmgmhMIWNOR4nKYp3mQnjS
AZYRoSbFg+9Z5scYNT1O2FPsHbmkEBdaTYSK0+3r+t6CYK3EPouvFH/hUsS6EnSdWV47vZJPBP9k
h/P/ppIh+IOrI/b5UkqjH+JGLWTU/Xak5I/3Oclzmn/YSjM8vx2N8Alv6x6/zJKyxPVf6h7PYRGZ
gkCTeTvF2A9gu2m6XUtdLZlHvIkVl0HLD2BSa0Qg6KesT1pXeaPFH04WE0AUNlzDUAx4Y8oRCoxn
LpscgltQbFvYPbrB9MTLzoS50r6JGtshcrBVpbLe8drbOgReS52WUxn5aCbumvQNc7Vqe3OMVEQM
EtAqLj76VhGFCJC3g6F+eGCBamUZAJ+5liFSeRZ1ciaZvj+QPoszNplY4iGysMXZttmze5no+d8F
LeQqsZOEDqo/gCqamwWs47xtpJZLoiYFKBHGK1ZCExV5+n5/eeAy46V8aRdGcHZXaLA4cyMRNonA
Kucnp7cxxB2eOuJf4I50K5+dyEPU48FYCdqtAA6fVbdzEcKJ7diG8yxbB5AjLMgQv/wpbQAAoG/u
un5hSElkSrE2O147VJukdRPuWEBs2TPJOk56yEltt2C5JdKN2REfuL1sZOr1dHSRLidSARR0303E
jodz53N/QQo6BbHIKpUzKZX1IunAV5WhDknl3Z3PAhRl1Mn6COfeaaUK2dS+4l6r52oQRziUMWG0
2i/xY8EVRIhE+nfSn/kYVxuV3gucHV+SoiSNqDMDeKc5PIOg9wtarpgj3fx6dynvaS9f4hh82rMp
Bvb77BfcqoTw/RAvGy8GWA68K1yaUPW12xE9aEokUfUEIFaQlAGOD8kr0kuQwiMSTNi98Bp6qO2B
hZbeqGcjgzlZ8SOqNdFRFLns62c0Skx/XLzhkUzlS3HkpSn/q2buhAdhU9omopR50fuCV6i5qI9r
wj7P5ulf++2ADVzU3GqpHjSFkMy97U/ej4RUormtKvqa/A8f6hTec+f0GLZOPiZlT1XLhkps8TER
tB3EHlmgJHHcxZ+hoEBFB5c6sExfFmvDHnvsi3ldTG+MTtRPXlMhqxcdj2QaQYwm+fTzJE711vzX
U2oXd1lrtlJdijSZzJcQv456OoOy5Hr6bZZQvZmQlDxvgADgN4JXiFv9Jum+4gAZwjHK317Zn3za
RK3CfZUOeuerlhcMb2A9tziAswDt7c9sj43wFQfBT+gD8gQE5PQGlctDQ8U2gU8PjbzxtXhda+Dq
yNOH5+d4shVNjHoAsA0CV+M462Ej7bcgzPG2s+07GVNDDBQNwi45pmDjQoV+MHp2dkg6gHMGFD83
nxseVZY2wYtD98aNdOqAQEH/lLB7M4DfoBEDkOfChGf+Sv2nG8npQNWrN7rD/f3XwSQIQYFiWaDn
76SuFYGVt9CQ7AQE+2KFwhlatlIwIONaZoPRqhBrG09LIhfX9z95SGXK94tJltgXnEyjtKdREknC
/qOkk7vzU9ExRAiI6RHOxTXa2qgAtKNSRCXqNePCytN97PIX62L0RNKKzjnLKGeKSOPzVgXRbGAY
V6rYYlQB9qqvKgh0Ncq9sHhJpVbzXBqvGku2+fo0DRE7ub5ZkawmXajEIpZ5fdkZtLNFHrX8M0MH
I18zpkiSyi/Ap0N2HEKa+hZRfO5GmdD566MTLs4x7mMRMObPoL9AohWo41wvyyQNvgk36Vq5weuA
rU2pGcGZZYkE1bAl2MxMES2kOji1DW4siTkDYXIntNWibnKLicvh/DK+tdnpDoPKVXlU7OA/w6JQ
nWmXH21fdvewzHjOqzl3W1vqjo/XtiGaLQe73m6Rn+pv4zxKRBs4eIp6mL8Sb9MhS/kX2M/4ifm1
pcZLvsCVJC3vYq3hwf/LOUeIG3fiD5aX5gVpI7hu+G5Br8WsM53txsh5Gp09fb9dKCVqeVDb3eja
3LO+mh/Wn6umyZuPdW0OACHoyaDrB3nKAGnd2xjBJZVzZdvsOtuQl37zYbXNF188K9yIRFVFwhPJ
hQ1tKYfD3nyJ8WkY4Pfz8XB+8/GRJc8E5l0cZ1gkXW8WpcnVLN8/CtmF3ReDYVVFdIzoaXpuPfxc
80QOuRVczWItS85V0jD7ZfQfaowKvNhiOm3lD+KgCzb8k91GQ/jYW0qvYMFaaai/X0TrSZDVJ8Oo
GwDKvDaFYDgMOGzyYTIxmYVZIOroEWC9Y8nf+JF9i2tCPZm+Hq+5uE2SxIs9/SsGEieANipVj0Bu
idQqm1KBIQ6bJvbxBfNHHs7VXTAFFxTFQpomxfPk+G9SEsAMFTKfGY8nncrbUnZfmMXDCoM2LVKc
D/iFXatneSxF89iBmqxQLDAky5t4U+AnKgm6w7LveylAXwyPZgNQeG8s4+Owi1IO+95RWHuqXKql
Kdz6sLWffl0FsXAAN75BSRPp+9FTTXeCqh6hY6ZtUWyswWeJ1jdOCK3B/yn6BqgQzp47WyRn6kK4
F62I9rS1YNrLBBtIwNwFHw08DQ88WkRFB6rptonhq75U5VrlCh9FUl9a5YA7Kslmb9stGcNnKr4c
KeiMZ2UzO56kA2zC3kW7dtBDzbWOJP1qngkyUrUDFFXgtvd8uXLgB1dqrHYBF1dgeksnjjmsQv7h
JL6oG3idjhaGmnQAS/OrmVvonFJSBtA7AMwUEw9IgtNVbyeoXwGSwqld9KIwmKLAx6oqEHLc8Htj
Emv2MAckHz73gUGnUZLc6PIYxUaJQ67V35SXzS2V+QF9bPJw7GldlwwazbK2iDzgU10IfDilds5l
CnYbYl1ykv9PzlHyRxDcup+vKMkLPhJV/HxDbmXA4pqKLpweJgPiaJ09mHIakJklm1W2P1heqmVZ
8MPs1cdsRWqzJR0P8ccbQ0+0L9Jd4CsU/rhu0zKtMyWC5XzsBNTPX6MzogFKfvHi5by77EMT+S3d
cUvWDU1rMQnXvzypVznWdhLbByZDr9pQrbqDlth/dMCDOAbaavDAUV7c30Nmm4D25LA8p3j2k0nA
tgSRiCZU1sDfsizi1injp1cpmAot2YuhS9gbk0RpW3fpylDnTde11Rr9pEvXbbVQ/ztB48TeVjB8
ZZBrmMdR8h/AmNtL2GAVikb/eS4C6pCfOqCoVolcy56lroqaN3yytiiLdAkwHpW1lMyfqgPy2wye
LWroZc/EchL9LPeSmVzlPxNfthYo+fjj7OiNWkRak9EMh+nXX/5L4WGsbh+Swssar4GpTwZhj1bO
c4ut5xh8wI/kQPHE65LKUiUBUXb/Mx03PRwr1zIfMj/2t4q0ZM9UOIzTvRDyeO8bYvt+rVusAal2
o234xf4Aaqd2bmI9S9nRSJ3Z5AGKC09KGDgXCFtChry3pHibYi5tJoA6E/owJpwqNVLBig/6ul4c
9ubY0lyI1p8WHmVjqijUYWWVQNBm6inbFqJYEU+sJ358/3xWnPrTc+5iQdHl6ma/8/7Ku63vYGwv
rejTMoKkgnjZ6V6lyd0uf6oX6iLu0d6g00OItF88FKFRWnhWNOrvCdJsHZWho0tU89w/H06Nmm+1
ZLgxwxKkGelCpCbvyNi7ECU4ZB9g2HkV+uiIWJVMVW0aeFboSHcwLGipAKxdolqrBqIPeKLMauQB
wfEWC+jn72AGw7StbGP6hZ44H9tWw7D7GhwLceUaxAc/A04ScyR6wMs/f74SECbjgzb1Z+Co2ta9
tVz3QtUsdMg4v6komy2Rlwq3bsV8IDW8klokhMgiW3DmrIFF4ePWmOF87R79boBvF3pq6VVKYPZo
eFYMV3WHztaRhe4zShRnU5YHQCRj6TUx0fpWtgfX1xOAfXKhOp7R6WhdbFvNMcv6EGr7/PVOJhbz
AkCkiaT2DnwxKwCT2rE/a1c0hrgsVH5LkLtwyxUcOU+HY5bIEmk7J49DMHdFlZpqEQ2GTyYjQ3yt
Lp5ZDSHB1rzhI87tLgzu4bHEktfMIRJlZ96DySXi6YdBDKTHhTOMyOvRO82F/V/qsFl0VXA+UvkX
lYSwJ3RDxxXslUSMqZhgs1zWGbgS/BzBJmy8kzptIgDMFeTBzlIqNkzYPDvAHR6D4M03PitsiCqx
Y9szWkyffItHDtc4gB7p9ZxlT58NlVF3nz1R1PCqY1doxHGCvnZkmLywjcgyP0/0cZZcR8up+GCB
xOb8CP6aNXhGLScVheA8PczsjFqPvfSCVKjpsgqWBQQJHpaoOHnvCusfiMCQNKeI6DV4P19vihYP
bsyuiUgI5injwSaubYXcXhUVNjxif78y39gjzLgCYbcbP2Z+cSpKSkML4b+julUMmFlbYoLLrDim
lxrOgNOuK6+N4aN4d9kjqwYs6VeZ2x65TuvQAYL/z1sSb6jcqVvgEajMo7rDd+vXa3vUEcsgLv84
+1Mp8M27oWVtPSPz9djWGTHuckRHBJRTqRWk9p6SO5TABWFOggDnYkLfMAXsULzadvFRaTN2Vu5p
kVxZ7oQ6fBDQk1X8LODxYHDax9a5XVtYovBpATHgpBxw9Ju3dwJthgOMCAxl/9CKLClMUOHqqPKt
sh2/020hIo/49aiwSe99MTQ/jgzFnyhiSwKlvXl1Hq0t62qAMDekjtWE1EO6PTriXzc7qtVADvON
Ti1j8veAfep3H2mwUVxq2g0DMvEGh+Qeu52CTn6wnjSExsV5r6flO0FXge3rFiYTuTiikUIVqGxx
FebutTigSpWP5BCb40tJmLoyNSYi8E72dOu7he9KM1jCXko8UnzLvYsoDN2hIxldsiYB95uOkeDA
E5imXyEWVm6haG3+1OvLNwm/MZwCXwcJHnZYxQdPKAYoaDSrWx27aUFJLW4WQwa8+/rbzNfLf/G+
mhrRH51oZ0sD8K7Fxuv7GYc1+tnoqd8+vQ9ycSd8l1KJUfq9ZhMb28krCTIPjrH2nDdrXhQYXTsC
piYMezpSLQlbS3RHGKdfNOlcz5DJ5HA0w547GRTwmfMh4zbZYChx+vhwnVk6l7p2J38+qYeG/yRx
cKPl6trl+4tMRRdbxDBy24e9vkeKHpEJ3NbB+Goa/34BZOWgfDeFHwVazy4mkaG7nzgChiii5jhR
KBluCTlhogjMU7A1Kl1SruKATXBhLBgMKxi2D8i4IR03P4+DxEYl/k710WoCJt50pX2fES9yCHhf
Vd9ghXDQl7DjvR++TMYHqgKH6gjDLCwsFec7gBspJ6HmdgyHBUnWbaYZylSvVRDzXvFybMs+1Cn9
qvnJIdGw0TXPA2NqhwwLPbOH2CNE/lSqbhbapCZOE8p2BHaWxr2BD7vT3Y1Ev3H8FLSg2akSNQW4
syN7ndCmVd7mitWpFRkKtd8DzizPaMyc0cjPbT2ncfiNCGL0SzKdxedXzU6XWV8I8Y+qUzw9qoF2
ziBubUZiS8ePsuwjcH9ZbwsT+WOUZyieDF2Tx30pYPeQDXOR2tM6rPu8I9lxalzLCMmy1N9ANljn
PbbjZFf25G1y6J2Z7jJ0h+o/FY0bc7dygiv3Lsa/D0/PHrRgkmC4HgP1VRoO22VYOLlqfsN2h0nl
n0Kyv7/DF14b+q5XbduQsEVEjJjAKbm3zcWSfw1gw0ZJRVykecVC6GWR2vS4ABvfYcGEAdpzxDve
HBpeHD3I8+MJh04TRyiQU2yvB85+XJ6mWcuR9i9T6yGwkerVGe3wpx5WDuki46Tb5v7uJmVUiQpC
VP9RRvDBYMkcENQ5TFAbo3C91JfKZ9tGNyFkabgokrx9hO2dGvDR90KyMLUAJ50myZe7TX/F4Unr
PcgJei29MPZACIcS8m4AzcOgcyTWiJtKc4LKLcK9U58N0wGCXhD9BvnMl0BGZlNiuYj6BoGKD1A/
0vkNK8/Nn7EcHlxidSMgvVVTeK4AdgdORUQbwECdHRKPf8BlCZ7qNX1um1qXJdODezT6O03chENi
H004uoPRu952qHeZaz7Vab56HYp9Ez2VUjNjoIVB0NbOSYe4OToFyutPASgUbYMxzf89difIcDM6
tVV9DW+x8VJn+PUQRHEZdHIYPgSQiWeFgcugo6oYdmwaOITQvtz2T0DE7urY1w/tnwP8td+//8NV
3cdsS+0A+CM0VDoPvuq55ZsWekI9P9TAs6q83EshN5oYNsApFazN+C4Qgvt4r4BMgOyyYAO8J/gc
Ij7N49YyCW+sFAaZWEcHHdrpcUMzYXO+/hHMNRQXSglERjX8IWA9Dx1ZluinWhaZujTCeCITJMqS
egTsYPvFh4EN5SbqDMzRNZQlDwIWC9j0s0c/wWJgYIfz/Sv34dVMXlSabnsslNsqN2fa2LO2rNDl
qjue9vFQqgD8mP6XHr0AHNMmXUBtY9d6zPCqIxnsBoPQn3UAwX1E0niBTz6IBVfHAylDssLsMEUY
QDKLeMnjt1wDKRT3ianFpOrEfsnIn04jqwvhYRsZ0ZC6Ew1WWWCiOrH9SgWPvP1wHXJOsRAB8HTW
sh2zAwt3W+SnlX9PufHJrlgwbOuq+IrQ9179N5KupBxAP8i2A9CiFX58N5M3jqmHt3qvWc9Y9KF3
Cp2JUI7CiH4RUht06d7jMwBjgPjr0rPYxRH3W33vc7TtDuy/BLjKpDr/RtRPY1aEMg65d81oqTo5
Wg5cFM+/8kV+NAxNf9gyvJDPrbw175a72+lrfIe2Vqcc9XfNF5MYh60itdclGbOJekFliqnWrT/x
+husJbbb9K/KlykXF4Z6sGz6PertAssfe7h7LnJZVOxAYPIqgYrLq2hCSmbnC2iNcBAhRCt3mS9d
zjZKtH3rZEfy09cZMjl/rXhbqj8I14TbK0rrV5u0ezUlc2wAsWdeCVuetbqdsQ8dr3CtSHLbjO/w
hf5XFVStJFDr5yxszM18yttG9TLOrAAehL7oUFviGsRuBnDp2HCM31ie76ogrom0LM6JBehKwyEV
Vmqd1eZ13BVrE1oBoSlqw6bhJyfCn63Cff9e/YVIkhWLhByTxeWV5xTgoPCLn+o+3f785xrPRnvo
G7jk50R+n5NBhN8NmazFm9WB29QBMaqq/buF03SnKi7JDn6Y4Ja0Nhe9PIBQiH88ep2JJkq3lJhB
Od5JY+eARPc5E/81BHxILlebQ+AaqqfpheQGTzFDVh4WFeaIZZ1R00PqDZY4zzliCxXselt4P1Ca
5379uytjaVR4B32LlE8VDOzxoOuuVr6/+4O9DkNKHJhgdwmXb54uSxE1d+HRuzRgBGAS5f/NVETY
l6ylMvfKahLehIQkAWmvzuhCXCcOWzFaqE2jwj4O/4x3iL94k6c/hlW6nKzJLQpPls0ye0Tc2AIP
TvVte/RmUsLBm+m/ock3BC84vgu/itfC5zY+kNXELyxE9MNqHlFBgdMDPJHOISOJciwqKi1xYQ1n
ww0nM4MKRaKOrX/9OvorYdnkSIWCmhABT5k4BHKmc+E2304yOFMIlp6edRDk6SOAf8mNjUkXPDFS
tRvNv48MGRdPPQec0VxRm56kY79vMnlCIC9B3nKVjGYVPO2Q+BG19FJdIfq6/TNvj80afdKq0zXY
4tlTdm8JgQ4Rugdeap3L+LzzYGd/5ae58cXZ9exAVYXVti2Mj33kZ8GN/ezyhIVUUadAB/HuPMDv
YFAUMZPnIvaAfKcix/TwVVQkprv4WYVzLIkCbvVY+nsT9eLNeVUlIQS/GTADf7iGNIi43nxgH/LD
jlZGf1adXAJAAChnHzkafA8HrpZaqSZr1gOuxwmpRgEUz3uAdeHms+j/uqnjY/pcr7zn+HQYfBmI
0McIeurSzk8ulhZcfl99A7qOu3E47pDUKuv3kyWrCsErZDmz27c/E546Gbbqv0PrrJpFpbooRghg
cfQ7nAokVi4mDrKPrAEq5/4iUL7HQOE+sStMJFUaeuqvlgPRdWBfqqMwZbkTpFtivFKuxPqB5QKU
I8BsM/ui7aXfMvC+SiWKCVkQkIfkUU2OYxZnlMAoPKw63wjcSLrDSAysrF4uIXLOU6zDNxesBPev
0dLAU/umVj/Bsa7It5LJnbQrKJV1SqYY73vIR0W0eFBW2CL2+KoTg0bjwe5TxZr0cnwZ1gEGkivP
cxPS+SNFDP/j/hzt6JZLEQAen4gTBYulITLDUVZ6fXzoYM1mpgWb7epvss1pGYg0AOMu42MIX04n
KfP6Jfr2JW0Z3VU9zdFwxyN/in4M/Q9OOwdvxhjsfo92c3oc7mUh/bjK1B3GoWGuRZ64dAT5OFny
LwxhDczyZOrYIrcCPqDy9LjYwOnOabwXvGO6S0gT8WS6ymBL+ExxMXFPqlNIH9hrQw4kVpDIpYPD
JpLB9mlgb01SzLJzHzNGDGtIYURxN7CZPlzDxMBnPNBtvrKwUvWIneR7ecmXkPxxKs6O6VS7S4EK
LzbNOdxfWxHSvXSNHLU1ZMttK9UBS3eXYRpyOvcv06HWDzPo0qGlYNThjO+BwJjYwZOzk9cecd37
ar7Jnj4MrG9dCD+xTpeokFP8U4yDaxG3C0gfGNRHQhuFJikqWPumNlg7NlLg93SGjoW7Db4imQDT
ZIi2RMyrtfDTZDrqhqTRVGeM9oEzLR1a6w/e6qAD1s0UItMlNGmEVEW3Pc3nycfjwFquxUs1hjne
ycxgBy5ZCjyyLupq4oiFXq6h/2J9q3WPt6Q0+WAECzbsfpp4LngBlyUs5zdAwbXcfNJP1O5UxNaT
8MLuMkB8bPtin0n/afGLZQfnJdr5dCcaMP77Kka+NQdteK6lMAQ22gl2DSuOxJtexjXiBJbejLiD
rDDzMp7PG4foXQV5em27Ud1yIL995TMOhgvyjStfv+/0dSIRB3iORltfcBsvarDegc1XX+AClHNy
AF19/C33Su+gwvJaF5NwNpcBMOwtm5YKOH0zMY795OrWCVp75zdnBBQ3slFuqt7FNGzVKsGe3+1H
ebB9YfwqpVKUm6rj9L+ddZk9y8pGb5A69HIiBqN1ypFXgTDbXrY0eG6nA5sCtj3te15fvhrqPEWZ
R+JV6cvltxzc2E8TiQ07U7iURk1lkIAI5AXDlH3ES29mdKixHROKq4+YH4bKjsgrGmjplkWvEhj4
ztVGHNBQXQS5O63Dj8wTuZhB4wbMFm8C5TL8BDUOjC2wWeT3AlogEgOunctLFFfAEzs9nKuqDyTe
0UeruuDli28o0Auj/LhSw3qcdIdHpifU4d9o7ztRp1v+2Ho77ou8Q9jbpnlFbwSMl1SMaT34Jxz5
34V0kCbdzXE+7Db66a94LtB8BofUtrOt5UdnyBsDYPWVxjtHh7T9QtdnhJ0G50pHWYouKDFs1WJq
JB8k1PImvurusYsSJQnvqRnTKHuiS5e+Kq7Zwaayelm0+7juzaDPZ6r4gi+iVO5T9qZTZcYBCNOf
z3xyYs5NOsx9fjsVY2ItdzC9cSWYdlMkW6h3ElyKzGuVJrFWhdNm/qi0LPOA9Rmo+ctMBUWYB8zf
fXbN6Oyy+uoPYnoiipbe1dmRw1zhn2lc3FU71jrLsj1V1Yvs0hypoSeBsaNvVQ++ERW4TqswB7lO
FhDgqmIzI7krhh4lqBOk+oZxNTMsZgLXPm2ujAKd5FlF75ubKH5T+B26oAETjRQ5nPZlZo/fiMlP
mFaj1lcMl5PVa3YSZTjzb8Plvep+2wX71E+4lO8j2hyqM35MG3iGIZA9WFtkVDrGFPYuo5wgJjGN
erBN6srZtXxoWvfi3MQZsPuBusTZ7s+fcGeb2gxNXDFuawL9nxDLumccpFiKayjpWS4i0GugFyHu
dcVKvaCk4SaXaVnIPU2TXV6XeuhJlQWIKu480HfLNFYjrVl4Ty4yM4+4PT9n5ItOHn3659mtcitD
X38F+zbq0kc+bj/2fJ5wv6Y0NmmS46C1Q1yJY1c5boX5iOA8o8Tl3n/TZ5vctGXJEIeVU+Ax7FOO
84ugd1ITCH3CF1nyY9YP5nAt53BiRG+lpHb0S/VAK5DMdiOYpZLtBsoKO+QMkdj21lHqdZCEw4pe
gjriWzpp7/VeiBfYNejQrv3OqLpQYF+vQGXNvAkyGQ7+ZDNedu6qcDQQSwR7Yk6dv4U19TR4V3Fr
4naxYY+AyVc2Drj3KWcDhFbWRwJxhT43FI0I/MaJ7sQV4xIFjWtMZqd6cfMx/6asbJWFJ9DEyaCs
sQO6xxTWP1RdxLAgGy4T6BQPdf1mmvV2+P2jrdDjvnmmpIQik8Msdy+PcpZJmbjcLSq0lM5/qPWe
p2g+twIYtkbgekyCKdUB6RZaqnH1ZcpbOplDHbG3ax4DpNnplyxNMB5wmdQH6G489b+AyKSkAKIP
g6xyNjWm3TuyOw1CPkpK9TISXpmJVTMVBiWF2Nn/KFeUyGJTYSALrXELCr6R4N6sPvZ7u2Z9ixMj
nZG6Y6wd2b1v5pqghCAFnz/DPTN1heFJ4VLG35r9VFmorDUAiMlPDx/Xec+0TQdU1BmwD7a/8f/h
X0AP7879SWYGelTxRLIQm8px4AolImY++2UMtqS7tgiMjObFAG+VJcYD/+pEu6eHlSjbdYa1mH+f
w+wPAO7QDfmkLo3+w3TA8eQf62ACoBE57zUe/b3yAeoaYvu4AW0xWkr7y6i0GAZbJ6r90LkM+EvV
BJ7o5N3NwXjPQV0RMBSqf0pDBfiY/UbpZX1tv1D9C3jz0sYjZOlAXbEhRrN3fB1/tOtLbWiiVffu
UHPd6rsN1znYzHeM+vUb0rbw9dv0FLmVn3+v85LxzTWy8YqcSexPH+Mf+c6glFt9W0x6JQD7qz0Z
seRnbnRj+WXICNgOJT1BOlzfvzLIni3CvV5bYvsSfHKcWw/o6HZhgQsEeMAHL7u77JYdYZuevICK
KDc7vkyzLhp54dpCiFGQ16PNsIaX4gJlbe1U1pDTCTpfD5pJhuT7tkXMYyTeKsVQ8hW8TgXA3Qbq
rGF4kg+q0ZB+1ZdbR7chY4ioa3CbQ/2H+9L/k7eMlvItya18medNbdcCGl/U6Izk47pBG59bLeEM
SB6N6d+JYrwQamVJdflmEdBIqrLuGlDh1QPRdlzKuCLEOgsv5rFSrtdAwwMuZTG5R/x66VsquLXY
9rB+TFYctOFatG+tRjkUMvewzG8rECEMLj5CQofP7aaRLImhCHob6DMOIZmZpUKScmCqZS6CcZdR
JgDVN8uTXedqjcVF1f59lhXVPwZChWb+klIL+5YL/SLUknF5YFSRjsX3oPSacJbb0l55o27lB+mu
dPtN8Wcaa8Ampe74+Tr58SbkwGZPhdBxdLET+Q0MX6G7B+fShvQqyq+puO8cOlewwCmqQg/ed94J
YwTlw7pDRlickhG6krdL1VoJuAvy3OpZWnmPEpK9OifHyB96Im4zCGsc+VQn3jhwDCNRFXglvK1c
hPslhEKMG2ytM+apsNt58k/BtnvWg7ErOd9aMZ4DnWUGnaFssdTa7U9cV1nTA++2EEQMt3pgNiFA
snfuZY1AzIyQGCkfQMcz/573eSjJ/nMn/oTG29BriMmgmKVx1ONQHGtiNe4bsU8nVR/WBXeeGZ2P
TgDxty3ydUIj7GU+lt2oI1p8797JFQWpnsZUTRMlWhN4W1PEdJF1f9RbeEjC3yTGZnMD9LSFRQEG
fjGai/rCojr8j1Bd5kiu2top+weevEwsvI9S18UigT/yEsOMNKsO4Q2dItBmVeh83jqvIsRrXPUI
gP3lYOwwyqUZ3Ge1/1P+haE4Rr/Sqp/kI1cwS48gPD3kz0JfNdwuxZZUTIDzJHj809HK6f31hP4e
i7LpjZ+L6srXtZ2ZlrCXLMN3k8uljThwGflZQDeRYEy58eHRYQxcccsDc1+gQoA7Ua5oWYgYPKIF
eL6sfvkHHAPIqRvWzC04WK0pgQTMNmc5TvUkmFOX3kHK2RcBkXtw96SCaJ4eamo1p/VIoPxJoUzG
py2yy1CNkM9H8hQdmZWyq2PhM+d0YQ9ZJBTHiTFaGYtUNnc7rKDpMKBvTSooigVWRUbTkkEwUCZs
LPKjZD9XZ6jb46mCPV+sz6/Yb/6FlooVzGSfiWY+xP2ks8W9sw4OIqq8k4VHsw4+U8wCJvJkm3sJ
WyvK6CjB7KjaWGg0vd4xFK+vfMSJOIEeehWag7fwdmkEAqc88Vexq8kikwHPBQnAZdgCXBcR2JhX
vBJqQsb5TvesIC/a7YkVqlBZBMU82CPvMoSL5crBdsdGkMLjmZwPbnL8nEg/s/cGn8cHF2SXq4e3
qk2URMFArsLvy2h6ti0CXEKlxDvmrsRDNULnMIqHwjz6XKAAyEf0s0LPomMw7ECyJ5gLF1Vl1BxD
aXNmnge+l41auGqKDSV4y2+vcoByI+Fq5m7FnA4vaNI2akIftKhNc2/9mpS5irKfQOpzdVXAS8tl
FxtokXiMNhZkMTil4Rl4M+v6LVZBCOpgleLoqh+blM9y/EEAisFn5knrljzzinhsjsYi2QT5N+Xr
Gy2vH5XXzNdc+DLVvRQhxu7r5aC1sQzD0IrLMDHufYHem3nrkpmtmZD01ugBXMrX/16s6QmgpvK9
aoWvjj/yp25tdzDxklZqW3Fr8NhmtI8D95cYt4gc3KCrrxv8uCThNAObDSOHe4gWGiVjrBsXvZMf
XPGssU/YYac+Pyt46Z348lq+X9w89Gx77uJQZDK3NuxVhza4ICW4/jjB5eLBT0IOzs33MoziMG52
UDTlUy77eGwyIDsCArwGuB22Cg/FzsOjDVeZoAENyYxZZ7L2Tj19XtBkkQKuEabI7HD8HPyRdftZ
cFBvixVObvpGZ4BgQWthqFdBO/ZyoCTHeYbmuA9jMCNNl2eQn1451qzmXrmwPZ4cQp6m5VgVOik2
JE4xEo+luHSXzSp+3gRjFmCsavxIc8xD3l2hf6tWbMqtLwosg6ihltB/Fw3T07zM3RhcducRYBtb
9ds28/ZrTDIusCXTMOO/OUpGvrtChqNqvz+GPe+/faMiuYmYUxoO3nRb0x848T0Jn6sQw1HV9i0w
Zu0qh9fA3mPtYq0uC2Zt5JF/6j6YhbSZGJX0oqICHH8GyQwXQPCmTXpVpmN+xmj9nupG5Vwahtag
z3N0KseSmi0K1keKQfBL9K+jFqGSXFVOOqd3bj9hGnZ6wIhy4mRGdJO+h5bjd8RttjesqX71Qwl/
DvqaVzp9ZqvXcpVXn3seZHII+fcxQYzdvXqfmWTFTk37aNc4xouBfderpjrftfcrM+1xNWetiYjX
v9TMW5iEQdjQRctMqh5Y4MwHRZD+KoYf5CphcPPUkgmSROzlYjvh2B4cPp7ns4Okld4mIRnQSbjx
NSJASkmTyrWhQ0b0q7aANOtYa1bOBd5VufEg1OeJ8uTSPMDPJmRtwkVggHbcJP7354LroQB5CsWt
LflCaaI+sSFQmHc1eOpuqLffDfbpdiAzCiLdcX79DufaqcJQWWlB2p8aDrZzC45q7JCIhaxSRLA5
RD8l99qWPmxxuKAa/8BVcERF5BLMhh/A70ERZn/fXsTTMQS0mXcPcIn6bVLTMyc/C+0DTyH53Bjg
Hy/mABV1ODWoajIUi3JJAPG5HcyB9Vka7Ek1Xwnu9Oyd5FSmTaVs/nT6dktXeQ3ucIHgrNMYidwV
od8t0RiS/67cu+gbHh0ukDPyMrU/hG3HEpIVAwFkJ9S3mxRkqgT+0YpWf3LZZWa8/hGDnleUdOS4
zvEeEUfNrHsHFLEhqFl54rYiaYt74ZmaUaNkZiXa1oGjhz1HRN5W/0zXRpuBKAfNI45woXf033QS
udiW3lExeVdcsBjGjRXJg927+Bix8cd02n6zZ80zviUH3l7PjyEbT9NKz1DcKmdFDsFwr5wO2MeL
0mNFqQJ+Waum1NsHF5YOrro/pFrvS+ONwhvRmZXC+w+1i0QymA2NZusvT5K9mCZj3WFzjlrgDlv3
5P5hdR6smTHfbisLVAY2RG4L0j/y+4mzue4VYQfXzvKlkditPu7wG/6IeeilcGuCS3bwchbUr8i8
UN6cQplG5bJGFi8fvJIZI1ljz55ZvXa1pBHL7eHU3VxBrjxINlAUN8aQkNstAhv91gjKnOZe1rjI
qrZg58RKnQceRby3y/iob1Q7/w5kCw0KgwMtxqI/idYVmcH88WjFdDlgBnXYrv4xWG05ZLc/bhh8
g4AHmxrRaM+YRtU1aDAM/YzBHuWYlkR4XiKs3UrRUBg2KEFKIRqLc8zWZe2g/urUEjHLz6GJEVcc
UPauJ8cH5DPl6HGnXAFOS7BB2P077I/PRv1RumABUr5Z6vkPMUtBRMM1G7G4igKJjWA0So2vSmJ9
60U/zTqW/0Filn6vitvyKzECaflGAUKfLVSz9r8YxipYdytBDHcBFfKQEWXO8niLUZkRovL2x7sC
diMrxgnYWKyY/eSJmi7O2ZUahPUeacYu5HkxLW6Eo80qMDke3CAObl2fW8DaX0UhIRv6BxYU2/We
aLY0QN4iUUGVRP533ehKNDB1OXfO/2zi1NWMaFkNnWwMaBXPbW5rnh09FmzmZCsV5WrwHzqDGvn9
Q77kNqWE59ifOhUW2Bjls/vfMetVGh1qzIxYM6PjJxn3OLhkC4vTgsf2of+6jGQxKH4bAlhEiJ1G
/wSqnQafP7U2q+oJ7MXc0vZd1c8O94lVz2L3XpS+qe0PezUJXo4tvOlVikWNPHq5PuLeGAbNWYrN
acl74z1CPKCUAEiIsXhPA+GjPd9k+K7eCnvcipR3I+nRa8s3vq4U0sEtBB/mFFltNfxcu4IQJ6CN
X/u7wQZJuk7k0i9pYVwGFuDcQDYdFGvroS3xsvY0d4MEE2RKs/QhyIbUaUizMsfgF+j3dE5HHXf/
IZzSiro8CL3bDRQeliEiUn7K36Q5rTsij5qvHhYYcJxiLY1TJ43IH2tBIUHGN1mzqIcv6uv/f6Fa
slXeuUK0PLoLnbTf7n9BpjsueOUT3DaJZLu1lLf16AmABGmvWKDx9uDqYVXMKv4eKFR6wafPa1WV
XxO1ANsczJIhfrY/1kPjN5IvVUsOkmfUoq7963Xxd2TQbjKNNbD7xSDr9wLvLP6gB7w1SUk6J/nM
tprEzrAB4Xpg7rJ97ynZ1GPb4NHfKqc79iylinZ/N1+macjJnmzuIN8BRm4jpp7aD7OksEPHpq7+
D39/dVZh4xR15qvhwV3mj2VnjYXn3gbyjTemTcZTXDLah0CPm3rbkycWxkuy7AcQHW28ErDtODdJ
QsVWqrMXi6XzhDcEEUGIlgS/uxI51NG4TCekeNeNGhnJ9sHKLrZnmbBvxz6F5SK4YNOyI+80nArV
UqvZT/k+8SzOdM9FNdNtGul+l/Mo+X43+pEPxYgj5BxK+/82FleiQ6dMx0UT01yIw461WfWgseK/
AlanjUtfZNRQmkHxWa7p9uCrLP67l2i/2mRNaNJEr4gmdfcApFGUU5iwvItJxEtKQOwHnsKLbRgy
vcMn3MtQEBQtXZ/z7MdEjSqfWuJPAmM8ukuhoFh7+RTZu0exYWOHFnGXM+7cuEZj/KgzJPRsygeA
OWQIqPxethPx61VP7L104ZJi4pkkTMoNGXvPkJ89ilXIpzyf9XYKh4zGjHqmoNdp1ols7bDXWuCb
IpJ83C3Wjm9t+qD4sM+NhYprm0N6a9NcTTymgIxaYGTvRbG2AfKlRFQvo3CXKkrYNPuCFZA3DbVp
Y0mUNLeHHwcOsWnJoNF4y34Q9gxdKKRlqSoPKUm2/mB9PszZA+kNimBfJlRDmXkQJe2Yk6sRJLBi
fcJokGL8cJGjiUTi8v9P2Vwam+4OzLXHublGSF3CRuUjDyl96u1NNXa0FBdpv21QXR50TfwgtJoF
ZKEIpiuVRg9+MdILE8ocgswVRRRF5p9OsSjoLQrWAk6BzTX9HajB6y4ySNk4x8aTs5V4Y3tXHlEL
ITXm/aWF59Mxl3KlZt9fJEMHg3dcRXZE9TKlQGGx1PAHPg2JfmcjOBHbDbN2XD1es7TVcEEJX3iy
JUFYGBNt0FQby5shBhFVA6guVhYwGk+0/aTQygm9ihPRhDVyY18HSs82tjiMpZM59eRSAW0BPkln
4CIjZ6n5mGZ+Na7brDGqLI7mokhE9EWHDjlBYEq5c+ulfwrWE08ecR9gE9gm5+Jz1VoBgZRroMZg
qKoBsQs03PoiyJO9pyj274C7dtQ6M0XbgNtlvZs7NiBoFPsvWgqMIdUuwshQ07Z7w7kInqd1Y6jX
/HdyC/0ry7yOsfNd/xoqrEkcgS8CMPCWHM8W54VIGjlVQ5fJ8La/OJy/7cHcXJa0MPO9XtRQ98mx
oEP9kAGKbG8iJfscOlXWVFClHONh9MZzvOlwkTVOKxqEHoCzTHtXO3fPQiK1VMW9FCerpa3c7Ofh
jKQQqRfk/J4U240xrxSE/5GkgGk54RVIRC7JbGDrAedOCJHzVaACIISTAXlevp21J5xynukdQ7j9
LfpFhy4LZfoPDwcPEu9l4v+cUBCPQyvoIY74mFOT9HWYkVskeFh/lZRmZJbtXAn/mhnBR6fZWNxA
pw19vXv4harcF6v1mgL6vm4HS/rJjTLQw8M17z2euf8Ls2mS7STgjDnk7tdrpunghyVjRLG3nrJA
kzmTM7tWPa95GKijhTyVMfeOOEyQumkFxS2CQoK3+dJazhZsSLl5zCEV/IaqpwDKTxPhggRyBJRz
+oZHh/jCqL6AoFJloTifH5F2P2yRBtVdTvVtvMqSM2BncaQLqPE6bCsWgpvHFpjCRlhSrvuCujFy
DOam6afh7xaKO+GBUbL3Akpr84c8W2W8noh/xMJnIBE+DXP01JD8pCj24DoCAst3CNLYBifivvmh
+cnIJP6vdEKULeY6JOt5BbeM+WLDiNfeo0xPDOs6xbt1XZJbiXSZUmZIiz+dwnE4L3UjAMwo+86c
pErt8kShrpzF1ajX9tWmq1sfMXv1mkRu2lzgpI3Inv2yDs6al4cIg3tJOzG0299SzT5XkMTBpZ1I
PncFXy9u0EKuwUDJkxbke5ew4cUmaNBDhuRCPbLDSxwMIo/6snt/gLqzRnpKk8OC/cx3XEHGONoc
e7bvgPeIBESexJD0yse3j1XE7NkMdhogLvca4VAjx22vI24lJvRLLZDpeCx1Uk/TawY39ejMydeK
5rM2wHX2HRC+yU0/y+N/fAcqvvgenuI+QTP6yl4fS3s2U2DhltFsXPU9wRxA/XTNGIl0Sg8Mukxf
s9qSppkG0zQ+OyXIxzhF6GTioVmiFc9s7qq8VQOovNn5W+xGY5LAyk+Mtum0pw3wSACW4up40YbW
CcDHBX9k4fwNvDaAT72RZfHXVj31xpmD+JY9WVLnwqjhK60M9tjIY2chq3h0pJVqQfsZ9MTibIas
G4nePzxJTQGCJtcd0vfJgbA0jYg7tOoaRJXNTbIJkfTB1dMNKj3dnWlMn8bVVrQUygMcMtlui5R7
whpL8MoKBPBbqgyNT9eAi0kad54/Lkw+dNUjK05pHjR2neh+UlWTOWmlFPIANUOaZSUZNp8KIcOX
Ptns17L2hdTuDz4o2X7BhblvOhcE0CKUUMoJHExkLlqjEcbg9tM0A2RUO/yqNjFBRXIByA+FlNX0
Ds5rW69u/WNg0j1yHMP4WHkmug3iP+fOk5sP2NvmHIPjeTfcKL+RlaFg9EGdia2Vdagj+XzwUiOb
JkUvaWPiCKM41R/qm/GnSI6qI8NwoHmGd3s2qPPAWVGds/KCWV26TGUKWcibYjQIz5ueOOZb0fKR
1MQElhnoI9ZLwREmjNQRHg32qWNZFRlgjwuPBUD8BYZmxmPIO3cwGXLghuXoZwrPRFpLpEv1ZRql
4Jtr3bT71UA8TrCEiZXUrVjAc855CqQbbe1iAwSSsuDxWvftzo0+wvvHDUsXqPfHD1nNsygHyqrn
4RzVHNV6/dHljkK7wD8Fj5U6+5tjXlB37KJVKz5TpNnBlWX0MikNwqatnfXlg9TNi4BtHp+FS276
YnAIA2Evadu1uFlpZGMltxAedGMtH8VT3DE0EGIHPG4cpOyru88DEl4YvNXkr00a5QgJTsztFohu
oI57tFLIf+eF3Ecf1VEHDV+z/Fegoo22P5IuoX/m1+5hzCqDoBYSO6rbRBqg0GKflDBLtScqx17b
jAFOf2O4QnKyEQmIFnDGurx+BhR8qzh53si/K8OzRcdhPqHnUxGOMxuZETyeR0ASH23/Nsw6T/R2
jVqZzVn2ytEU+GALXqDPdOMo4IMuxvXny6KOBbZOAl2eBlYPoXjg91rdqszEqT7FUOHwe6NIyct+
PEoPX9vtS+In5mOaNl/iRRYksnuc2fKbp+BQC8Tl7ZFXdiB+xT7K6K164SKIWOYK/hRJ1f8Yn3Cq
6JKG6DVIbU1RhjL9M+cU/9AmGIy5cfsD1X7x2Q2LTNy8ODXD4JEZsY981XZJ3Rj8LaD0SXs9RMtz
yZ5Okkd5V6UvptEsyfjUjwsCqjb/H1vpKG4nhO6Gl7O8AU2V4s4h2oV5FjvL0eGfCn8dE1rJFpXy
Sw6lCfPnjozBlY+Qz8HKr8DLJuHZx3OPdB3WXDU6YoGCx4tX9ipMxwe1xhWaUe12sr36O7sv2Gsr
Ko6fcrer3wM3T9bgHN22j04WoHxv7FME8/jIPNBJeWkuSZEvC3HpqfbGp18MdrjVnTC8+CGk/IKp
GN58XJ9RFoeu7tCB3OnbuAVI2eyYyg/1jn5ZE+qmoyE8ckT23i8bgrDlW8VbP+/aaFVcHXmFnTke
hpWeGGYglgFujz8t/AqUCAf7th1zpEk2Tx26tafPq0bxPhn9rxVjoZVfV8DYp6KFVxaU0823QGHr
XHSJHwxFCXx5ChGt5NcJ0FFbQRF+cIRHw8Zm8uCeTuiPqTP1cinhS3/LQ0LfpuuT2pgXHoUR42fI
wPpeVo9pvtk07fFMSyho8UKKaOEWZ97F5BuTlSgktTuZyp9IFK5gHHzOTgLj5LIt50Uzfu7UVn2H
HQ5MzgSXIkUVtJ19bl+8WMdXiZR3ycev2WTHAYdLyF8jPIG6RMytoBnCdRE1kLJYnCXKQT6Witt+
OgnC5UvWLZV+clWK0b90sWGeDEFPDpNqu4unuEn2axPLCbgj+K9uDMh7NFNn4rqZbk6zrJKiWRLv
mAojvDA1JaU/zVWoooFiXUlN3utqZjWjrAf1i/FsO5upsz7FWm6BAq5ciFzAv9BZriuJPzFcY+/P
XE9WoQ0PwkkYkFBOwn15v/yGBRlxxJqrQjd5yqmq73UOQbkP4KLpHR2vNxKKEPZz3nDUxPV0Uurp
rgaQOmDU+5/RCzKwKZ0WBpStqxGETYFo9/hnIYMcErEMjJhkxjV6cJcLXnxsZ72i/QiQvwTM7Grb
4H0oJSdyzrXVwOom8WLucKWfez9l1hnH7xtKBark0Jyfkz+mQaA//Rc640k8QwxXjeqqWhmjBMSn
502uswOl17bD3SI70k44SGxsG/q7zX6EwUed8TdE5myogssopkgzgVxQIdOLrgoK9RFe3p/N/ZqJ
RcTp+xe290Ak7VAFVr4ygLSeVHpjUUR46B6QuukRci2cw6aQCWeZ5CBfoS5Siz92fIxWjLNfzSUY
wvHzViNkuwNW8FClLXQ5F4OJhEdeW0YarcCB3H7BE14BR7nBu3/ExbLjn96PZfi1EupLi8ozhp1f
fgHaT9ZzZ5aXs/bc8GEILIpHizRhYrydHpS0csAXMHV79Ff9FNwi8f1A4x3b0N6xOsdpwyE22P4P
iwnEoxttae5oNcj8Smz9g0Gxa0iGSyHEudxeBnmKxapCj4YMuG5AqNs/Eosy5icZ0VocF68Tv4JR
fRSq0cho6RYrROIzw5G7P4C5e1Y+lMt1RMkoKcyzzka1wdKyMvABERmL7wQbzoTbzu5qqnipUcyR
dDjIIA0N0mPdtF4PlcH7ov/FE+Mf5tWrBHlilsWONM6mPl14n6nc/Zwf3cawxSv0m6mFg88kie9A
cBlNxqA8x5iaGY6xPVFywjxkZxhA2TK56ysxg+LeACjNnCKBy+DTz1lFlOvolp7SG2a3H86uMZ7G
UVf+k/kPSPk0MJCDoURjMjl5G9OIDMATupWo8c1nXncTAkD/0BLCXolcRvjgzraZK33hfDxf2vxB
Fxx3mtvqsqHJXuf1PAU0Oky3eOJi33i/NijUbG/6iQmCsbBfS1FIx5CbRlUsyqFQVDNZLJt1AWg7
8YDGdAxo1Hltd87ev3be4YqqcFibUYfSbHNPUmei7gVTGUuUDktxDW8mbCLWt1Y/sTw6lHHWTYgJ
9ZNZtMGxFzwYS/yg6SBGtE7giMc3UKy8BOXPbEC8ow66e2tSfB5ksPIqHeRsCrQ0Eb5Jm5OL6+de
j0RE/1BrJ7UjahDWfSBL4O7T9tkEOU2ViRig+ERZbdjWoV0dINXa5+YJWLrZDwKVeaiHLPmOPHJR
IvhZndFTY0w3JCvZgHWtrAYmLtqWyegSnT19hjbJD/NbWavG13Ogrs8UfrORFcwxl49U+Y389odh
OehZtDwqzkL1kUU3jJJmJOTOPCffktugyPmwPC/J49BrQa0uBFhoMJjJPEjxCbxZGOF1lalFE0RY
HqdxWGePDXhY4ywXjfCN9B37cQ6lpgX4lis5PNk4UHWjlw624HxPFl3+mrO/W//f5lX/6xqvZjLG
bL1JVGLZRaYdilVyk3ShIaU591L/PlWM8nGmX1sWyTqHG4rc4gnYkftiEqD76SzJhv7X5PgI1Fj2
oxS/LRhxf15MOKjGbVGNSiXoWaAH9n/pRSyYEhP7pBUx5ZKMpTDkhXJq2DAG9bdZvQDhjGDY0I9f
JxskVF8UP/4DzMBZL3OTiIvbTqFsVsSJkl5Pdfb+7oCZEubbzbJR70b4sZ0kSs3VbQdJ5Y/91pYQ
P7MpICLeqLi//1zBmrGDKMDP3hWogtAMdgFmzCYTTt1VMx/TeEv0nP5ZW9+f55S6X+1sBEAibWUQ
Xy1+rYytuqDpG3katZXSGEl5NweQYboafA7rKf6zT+sqw16ukbB0Sf/LO+C6/rYv73DIvpKa8o2K
kih0NBdZDCbH8sz0WHu2F3jTXWaOKk+L3ODBbBOrUq6HEwwJM9KR7RvjamyoaFdoRrIinzRtXfat
DRfb4KeI3qErIvNeK4aaetRmc2rRATp8o4mH9ELjnGH6Y917bbSIlhyGZF+3lf7Pc0KcggZN5wug
I9l6H//hfAw4z1tCX2SX0eAQrhaLdUww18SF+db1vCeu4Z5+8frlmNfl2yFx0JFIAT75yrQ3/RPV
6Idcp1ufO2MGsScbCpDeA+Gk4z6MZQFlnzx4RvuhDw4uHGb1LAWgl043dK8SmeYLNuGR8EBl9nyz
5qaiRzBHtRIkPyL0wfS+DBPoSjdkF4GxlEi/bCojO/lBe0i0jNIFZMDQcDb08ztIyxNv4yJmE5vX
rnfQuVrvz7IHSWdMB16PqhfWPHhOaIQn6LRnbQ4bP7VOe6wHGQa29OQ3axn9nHL1K3dG2BytDKMH
1zDzq7mRNBfuAn2djtCSuQQ6u/VhWoISEH+4YHW2lnAipi0BIQ/Jx/k9TopDPFXSnOkMcCX39tm1
pbLkWLX5/FsGokO8uMe+1AuwjBJ0nRJ3DJPNIacMEgVeOrs32qPg4HC9Q05sUGryg2ngR3G8Yukm
ENomF0xj+RvmXe49KpKvnEGs7L64IAZABFNxOgwSWdp2tIqy6k3rxnWX0Cwy0sC7v8Tt7f8aOYAJ
K0ZrBddf0RYDyoUz/aFXdOfgxIoZxuS0+cNuqChjTZix4jC0Yc6/XPN/zwv1jJdkiutXc9pHvuA9
DXe93vLA3nFvQjg16A58MG5BVyzhZyl8TTwYj3ACvFPgwyjP9ZyZRx5mxDycfMU7UNK4iNpj5pwI
Fl+EqL3+hWxzTTbs2OGlA4J2LFjv1rHpG+zzBsDLlDamzoNnuzG/5gLs8QW0/ui7PPxDtUEXvhKO
hBUv8bkqRY4gVXVfaBN7JONc7IBBF26AgJuFFFKrnyIpCWhGX8mLKrdOXpU75gdoiSJqMdzyp7ZM
YACDDLoqeY/bL3/fScwWWOQpmyx7E+KVWEFAIYvIqMkOyJ43tUrMdL3vDKCRvUZ0PytpPJ/+mwLO
AoJD1ssKNECFwDPnMPO/P8jDd7XYZjXzQV3+r6nKXewzpqP0EbK6tF8UW5j4TzTr6qN31BNPiWBx
NRPGryjV6zPGgHkh/thCQm62+X/9s2c0XaJP6gtseGP7H6ErVDLimrPcPkL/VwmhQ6P3HVOLDYgB
K29+9RY5KIMYdwuW+24JTjG1jD7cXf6R91f3naA/cW/QNeQ1VIv8p5hGaJ8CAqF7HioF71Fe4q6n
qZStV8zjQf/MYoEWLCDMKXcRxKsBAGM0va06/YRE8j+UgK+V+QOCVw5HT1mXr3sJK377ZzAqMeLS
M7AelsS+zpgTtYbt5hmrO+cWkmPbFSyYvByMYFuu8fyAeRTayGjX0CJgTOooU3BO15OJfciEfZBc
sqRFyqqqghmR4MqlFJpSSv2+cUkoC+bNS/pBBKCt+NYNUO9mReb/U/vIkbUR1lg3lmpoQt1zt5Po
H+Z9tnW2F/ab7FXVfx1KSM8dGjkErWaSpIQ5KyKhCChoFnpM0r+5qUiqQ+Kxz8d2xHV8tgMYpkHb
znv9eyIaQyVb6UhqUHFuY3gLcryKkk8olHbJ1KWx50vTV/Js0i0LVOZuVLViB0R/TXQfd2n73IkN
AbKGaecDIHWPxTdKL0c/fj4aKqK1RiZDv3l4KrsrMIfG4YINO3xSpoUB/QVTTp/6GcWub03yXnKJ
uWO3LDTXQycI2eUQcv+/ts63cUpnCJ6CZIZWUBqIlo7QfM3MUt10e3vRpjLycVdUnnr+l5wj/yeq
R9qDdk+1CxXhTmktidyrvnj6mSByX/2ky+UFbWYHsnv1wgbLP9Zl/z7jj1/95cFIAtapBfIm1QPb
qCUd66e2g4d0Q7Dyr/5iSSUvWdVXebE3FhsrEaffdcYmdUzmu4PAKbokUycJiR53mcnpVAmFex9M
VYz3LLXmhimpYy+rmFaGfpNt5fzzdHi0ket8taLwP5XM4G93QNuZuCUcXQI3OY7O9vBBtWurfH4O
EWUunEMedl8GmDH//YSMrxHHuCTTx6zSIv0q9fs1d4HrORoLfdnYtpmJz5oSwBOBY3V+StsE8gHo
DPcF21aGw3pylU455Z4YS6VLQIrpRcdr251QABtmnz9sZg73LOWhGeyv21+GmGl8aiCzOmcrraIG
7edHFX3leWlUe+MRc5SLVZaRk0kauQnJrQzyXasVncX1Ih+7m5GornM4c1EtkjN/bq/Qj92kXfw+
I+lGv8OUDO66yr9NyMxRXjex6234sWdrtoH3eWMiJ/O3k8iRyaLwB4EL3GcbYoHlyLS9XJ72+7g9
FN7JXK60oJmaSfXpk+jZKZG1i+uHuTdHhFbzVUgpUYuXN6B9qRmvc6F/s1wm3jO8FVjfy3xBJ5cI
HxQrw8X4Aq/QHF4m21FRi1vYwXygITcBPbCR5blTMEJykLqzayB5yswY55l5HMOsyt3sNAXKbUJC
SjSu8M/ZhGyfA8L6JIn9ga0wJb2FKrWwDJslWqUiIUf/rIi9wtu8v//CIEb84QedPPPzQILnQs9K
cZOhIE+ibZUeVnQUESF2bdGxnUBTWerHb2nwYyYwMFOoSL9ylMifxQRnnzEi22FRfpdjXI35W3sb
w/6L21Z9e5hj5fDCKz6RAvMN6NwAB6OiBPPF8xZMLcTdD7f7Sg2d+sLMblQqdP/KCDKFdwjsVpqX
rTWXavVPxnfTbsYuPm7U+0Mj8z0qtGrbR1W3TqBK07ZnRhHTjdcte+BV09ZEcUpkE5awr/bOQmW5
+E5Mllj0c90fxOU47iZc7fZGcbUggNDEwYonP9I6Bz38Khk5N8GRvf8CaPpVECpvSmN0MShQlJ4i
4ZiNftu43xHI3CPbFUeo+on1XbRmTd2Nt+dmTUXGRLfVw8S6Fk4Tx0U3oBYVs9grp8PuPrzp0lMv
E+jRyJ3kDeiQHhzOnwz8E+zcsXYZM2HERupcrnMHYBWoQDnKrz5thGsg59BmSJBZtrQX3laSqKXP
ofW+T/6L6Ob8J4dTivRnLAiF26F/TqCM0eWAVbKU5dYNhWIBL4VuITtUrVMLpT8jta5ELecHFsrA
t/0EYaG3Ysm2bE3vv9UeQgGGkHMP9mN4BASRazXlljBsJ8kNdDSHER9JXiVlELvw2ULBZZN9xMEd
AXHGUsVITT7nFxAv1UlgFzKPr6AuzAgOOwn7iT0j5NFHTMfSp+QTzD0jS6R7p6RKeceKgvOdedbe
MR1SKqJjA0PR3rd0O57D002DSZmP0PAP6sGCHctbpYzGp7WkfLbnQeIOmll7I7fxjtBVHNpJVw7P
WQ1p6h7Oo4VXFiQVMSNzVb8NTtnfvL4h3Jv88tuuf5IaKb802D9QSDPWfhwxoU8hmMjqco4KYL1K
ECBJWYQdGQ8Zv7yX7oZjrutfBj0T6PzJ4bRXT1bSFaMXBgpuiIuLCtvzBVkDWkxtUEfKklz9J2w7
kook4+tTMVgMwCYkkXqQZOqjh2W0j92bDZNMipdU1KX0u5iC2sk4Ro6CBD56mM26aaIFMR6PLsPJ
2D0fLgaegg1P47JkZ9jgownFO0LxZfCbmvkIlulsrE7YzjViyLRn0KwN44M77kOvOTphEwhS+j0j
61QA7AoudoWbjyZFETbjCIuHnmzyNIYkxeln4pSvFSZJ5prjG5LGXjPlaqQxaibvDuzxhmwW1IEP
3eEq//VZ0iZJZkZctiRjnj+r4LByZkdkaTnpAYf1pn6hSe4emEJ6haJXMAr2aAcIUuMCZ+hFwOha
ukEl4/xaV+Fb419nsnK2BqpBxwu9pCrf/+CNi6VKlm+CqedlejTaJuzkrB27lNhmF0/5TDQlQWxE
pOTuXJyAVi0b3aUf9JOFBR7+IxC19xKhYqDZH2IlQnLANwzBv6oy4YBVX4jnvUnt94gkgQTgbZFv
VGPRDsV+h6tquND7SPr8S8Lf5kEw6t+iCZkvlO/ipRg348gRUsXF02QFGfeLul3yGWmeITHjYpPF
3OoVTOVjXpvNrtUGPRM+ebowrW8X9FHeAUGRpm7UmNk7jAMnnZL+sCmV2DkhzXu5AQWqj1kWHtks
0cjtjKbC5kF2GZexw9D9G3rYShUowsISZi/SzKcAhKNaipnYqOXLvjpGuis0SDaq5NIcALthG3wU
XBXZRitydBxBeD5zOq+NN9gqCELEPqIaoJiTs70uZimSLS2cySgtCiaR/DMSLElbdskJ6gw/Jzny
fii5wolf6WLLwWkwoalZLtoZnvjQnw0EH5c5+WeK5eYe3rA2lSm2Gu+82Zke/DHH9aJYewuZeilg
s4kQqLyqFvZ9SfNDEueKcHeaY7eWDN4frXuEjrGlP/pzXrO5Cub6/wAUsTORPNTsRFzWSDJioqpm
ZaOaN30fjMtUIGbyAYqIjp2wob5eDXxiAz0RQcmNMN8VdESl09R66afv5nhoOQdckAFrZLwMYjQv
sjCTKd8nO/9yhJo8DwO5wSiPT0QYmt+C1fMSG5muLhD4t/5V9+OFu+fZ2mKEVgpiOuLHxQf00iWv
ab5ukPb06jzwVV2FvyJZryGjL7P1xzU8DP5v8gR0u0/8dykrVvxm2ztcigjVJyQFt4JcFZ9dq4YG
khC7rczZ0lAGUq8zRSdLsGo6Hnh9twPwYWKB8MfwrQmAv4Xf/VISNuBt73LvudvUUCWSoNlAMjnS
udm4lQilhdy7KMqBzTeWgKIKSR8PNwLIC58layUO2FX/A4amCmItVDQtP+FZ1FMaewX5f9ebtOsz
n3ufrYGWHd9R8EI3QK9iB5/8XHi+tnMt0dnu6cLKLfe9LFZceNh5hiApkQ7IMkXECgoMexOTMdTC
QusKblpuNqpBcvHqK9R7y+2HUDp9Fe6+pE8JjTV1JnPjGpeWordI/m8dRRRBv4I7R0fKFJTSZmWk
y4V+/dPLhIGWJ9kxo6JN5qny1BWCxZ+mJHXcFFKChRLMOmDCJ19UDSVCoYlz52ECC8FYXqFGLkBS
OltIYzSZlVePUuZKxLZgULQdL6yBcJpdPSJmxEvOOLmOdIWnvF38YSnYDf14zMtFw3xPLu4Uu6O6
cA8NHu7mYIBGwzxwHleh3TTsJ64qnn2JY3nBUHmpTJ+JtiQLcFaee704j7ISpypQBacHC4bOCtbm
wHnttyqBWUc7qcHEzIsrUk25VMNL+g1njg4TGn5ZtEWxY6mMOElw4Gz0f9LseWzAlWwC32yQC7FC
4DdHxGMCIlk0NcnvnKZvM5DvrP8cvDHNzD+GmNz2YyPmnZ/dklOFrtdbgNj5yH2+7onV4nTdDAcz
kkrJZFt8UM9ezFGZBCKXRT8NwuwMD/co8cuW8FmMrgie5hRg6iAI81sa56DfedrPSEc+sL2cUQkc
JYyAV/s5T+5mAdN4y1SkK3JmYZOO69e0LD/7SsxP/k5iLAL7ML1OUQASQHhUPdUPfLi6KGMDVTGm
xFb6yGru3knVlTaJrVqsOoeEb5g7eH9p6ocoghs9HCBcIksQ+Mu/9FuuSzr4LP13JuVBXA8Dp5rC
HiMDwMEgyqcfKBtyRvo5Jtnk24GYIMkAmQirV6+R8Fc4VWDruMWawFGnz91x68wDj5sjxR/3OCdd
GWzznOph8fyk4r07ze2EVn4fDwjNgLwpOPBsjh8Kwt3Vvhu0ut2qsf8t4na7/gCLF1nKjFiRXb+C
BTaZXJLnheY/dLby4Hx7U/p3MFDKYpeaIveYP+k0nRt3jQ0qjVnloY+OeLR73US99ivpe9L9eP5q
T0KYt/YWfwaSVQHvM8G1u5iPcHOgAEXzKe+vXYxHZVyXIpiXeRPTvbPgWWhxWhBz+xCA3llIrU30
1OXYFSCHXCCroAkwGaJAKKox0ye/1XoJuuMf7V6f2gRSRUQ5egtuBZ5+z09GtK2rx/jUjZKR4BqR
WWicujGMBg0yBpzBA0XsYUThDy15Vv9//IUaz1m1kCKfkP079tjLdRXbO2MFlZu0V4K4eB1WaSEf
O4JJ7PJXrpAP9Z6A0oh2vlBGKUtb5z8DFhFidvGQrvQZwl6rAscM5Km73KkivL6vn23IJVpWU8V2
ZbYIjrkhq1Cs80H1f/fE9WncC40VlKLWB8hwNK610sS1ZLFxMxFIQqv34lOBBfwpfn2oNNEDC+qo
vjddxjA9FZ+1dt1yQJrTlJNZFh5v3qifo9+B3xtzAxKxolryRFrHk0WTUDb7Q/LZk9i57aK4+N+Q
9oUM+2iQx5SdMUkCRY3ErsYQ2eot6Sq2bL0xo/AfJDBEz/YaSd3FkJa4paleTLGpmOJbl/x843sM
fNGLm9WW1ijrGXRxIJaC1lQi796wYymVWD7Uz1uIT7onM00LRy7tft06gHZMl37dfGrBPbedf0V9
0ztsD3BwlEnpyT578GbysZNlvRQjUH8MJNEzNNkSstuM5r0nKbynJ3tGW/hwwD7Id8udaG99ksNi
EVMsbIP/hDndac6Yyt+L9Wt6savpnGxqs4GpNVu2VN+k71hJPTQ0vgSYL3zIEOT91LRv9YIA2WiU
87hseCIt0/4VaYyfccD8Jq0JkFENdZyjSfiRaRnmj3gqJJeq43SqvY7nLMAJwuF94lwAm/WEcVTk
c053TBnONAesmwZ0TvN1G33RFKiAChAl2SVdV0c0oRe67nbfpDKJf1+KFMKhj6qoZaKHZsRou96p
jNEDi0qIuYZHVlsPLCZG+FrN6qUNBToTiBWFdyRV+YbOZ8yJSXKzwOALh0orc2K5RJVxQA4OfHjT
idEiJnAPEPN/6KqfBr6tLqTXZGjgyJZopVn2n4/S38ZaPDpHijBMu3xkm2T/tBjhgMeWSnpmoRm5
wpuTTA2SKrp3m1oiMeg92z6VfEcLQ9HVG8I3dtbyWVxog1vuCvE/RBDJZNiCssUTcaRIER4v8BBj
Ll+732SyXoF0zarvbKZBn64ij1glkdoW+mxKL/XT4Bs2klZ3NVlNBYE9qPj3fmRVwcB9UL0ZLwGS
BDONkIjps5SjQNx4PMkdBdOwRvSG00tI9nMbnld4v1MxpbqSAQqu5bfGUNX7gp5QoTVWu78HXzGq
phiGn9VLGfTzM8qqoUkDqq9lGWl9cQPmCmnsw6UlfpvKxzQIsrZK83ia4Qp80f4Sj4QOTpZARouV
Cc1TWgUEf8DjcfOa3X0Q0efh0RWQ32oCOQ3qzYvtlmy+3YBJv4ZMO7Y8oc5vpzvu4xiRx5qvBDsg
aWwsqPqWNCp+O69fCMUYCY12SGGvEW6Z4AARA1txCw5FxWhB1edWRX5uVM/uKGqrZKcl5z0wpE0n
iDs6s6Fp7uCV3VhqWt66O9D2v4ZV+6s2aTOMeNyFZ/s8LyYrICbtmjXLEtddHakD5L162+TNQuAE
jaDmnqjjvcPTXenI18KhreiyX5q0H22lapksMN0w/nY/DRWXrKuYG64bVjocIOmQK/xfVzGK0HoP
sdwHtbApI6Ex104evvlJec7fkTmvzVecZPhOfJw23Gbh14lgBadnZ4FXY/EaST4v4KE2uWu8G/wy
q7bzU1v4l/z9of9mtHcsl5R1rNNFDpgb6qTbTiD5D7fR997nkTcABu6o2TMAdMjSqAvdxGSNwYTt
ZPyUtbfqnZmbyDMUwaKqdFG3f+wnMDfP2oHrd8jvcVuWMULlD9VdoL1hFf0jWbyO8wxy7u9QaO9T
DNj8L4zSIGFpbSdptJWclbsJA26nywxKB9Kvj5deYyxO/ahCxGFehU8Iak+fXc/K/42RtFMeFGBc
fetAXrOWeeuPat4MaJuHVLNJjweeMJtEXZC8HE7hCo74q8mwYT+MIy1juSYmTUFjZTwZPTfDq1z/
6p3J4qcEnoh5jtbHWrpKksSnsseylNpXDgF/8oEJZm+2lPCFE6mevdS7uPiIuO7sGF12CVd5AsaB
RbuyGlBxpgfupGTYwVZiosLmOQECnBeieD0ltO8kEIZMirU0J3/oT+9L1AND+u2E80/5kPUFxTI9
y64HqOsodwI89O8OJD6xFIXojK7bvQbXvmPPuVRpl1R12Yh69YMPZBqornrM2Fq8YlQuzTaWS5wl
viI+F/7/ThCGbWaHbv1HCi2rp0hZwPqvtPgk6Hf8Pthj2xUY3vqtkr2cieuQ3VZTzp6d6lvPEAO2
r1AdLHrpJ7fOyO4Ej+kKI0gy4QQJaBVqAN3FwyLQB7QgyuY4esZGV4Lfr/F/4KBKEU1VDQtThI1W
oQ/NkBIbALfiejkWtLXHPVHovMuLeGToKhWEfWYAchsFFka2Jam41h2qifvQYRilmD+oQFVKbBWA
3rm58dfou78NELtg38fS24DxEpTFkIqpeC2vddnkP5diW3MzFF7C+/hVnVMM28FM+DTlrgpilBfJ
96k3FxZPp8WCbtkf2VbjRnp7CBSxQn1q1Bl01/fQH+NPAu/L5pqXniNsFpPI3w24Ux6Jgg9vmIoC
/JveotoyqR9fhJVEN3/vBPI4QU9F46NOb3RxLa5i+VOAaltBOTU+FE5NgcjtYOsPxtCcvdmFf2rS
8cEZNzJIbhiMMRj1PJ5/6FSnNYRDLmKTaZcbwjEaTyO4eJbQa0A5wy3BTPn8xz+4+BbWlyqXIt/R
4nAVWUBOUTnehXSxJV8DBlXEnX7fB7MGPn4Zd3hTr3n422//nea3zDyl0EaKHwOybMBUF/CU7reO
FoVLTYrbn0+uYN0zw29mQjuOmCic0GpgKQf934CoHtxzkJWLl8wjewSMhO/snP1CDAjfI0XHFhfM
KkBeWAlHit8wYY+tXXwQqnUeawBRTqvvRkZkcquhRuLqwY4m49GIABOii1uPztCUBNcbbvyVyGtj
JXAJvy6Rt8wgT5TKYmlWqwuB4f0lOLa45Zo9F+UVjOWh6ejtu6dXpqeUy6y2LFJnQZXE09ALfsWc
2YYE6fbmbDf9sMMq6XRqrITgZoni6u/LUjrvHuDlcG8mZ+PuDqjzTVf/wRd00hF3TMRij43r3Rfx
nFIF/DXWc7zHZsinchHT8+TbOL80vNWQAGV+2oW66SkbLJSBwdsbUpf3Adqns82SMJq5rE4sx+b9
P3dobtwKnOk1drth0ZzKEKShMzG1BNcZnyumzR4MwsR4lZD7gb7qL9FZ4xyRjNTaqsGYKLjYPKqy
egANn5A8HCImOyis4uy53k9gf24SB1xBL1QVHB3eQfg5N5VX0lASGyyZld0PSPxr3oE8dcdgtCY4
M5YQtrgqyE3bUJH11/zDNotFFU/ZqRbfyDD8gL2TamgIdlM7OVM+9XGp0Ga6MBkq7HdiYZlPWmNz
YgcXE07rPoDCFjrIx0q6S7BL9P9sw1fSEdaSv5n3jEnF+dVcXFxyRwcAkpnfxX0FxKd4P7H+aSsj
eDvO5/mEHhgjeAl1gIUgKq94qWwG74nzx1PcWDYqMX4M3gGG619BFa3GdS3iEHMGZyQHC7Qz7hlj
caEQ1EgqYOu7q9PQGqTo6gNqHLsxRftEIYbCtcsoSJ8eOlJzDF3E+txwzac/rYu9XJKVT+JsFKfW
ijr9gYJh5hh3c3VZQrj8Hc5RPV862/zFyqkdwf7GtOZzV3ZKpgacKA+53kKjUF/IBUwkI/vRwtUo
6Gm9taKJ0YrTu1bbQgHTg2aFLMuClAroziJl8AcjbQIK8gNRn3AeNGqtojlrmLYb2uhTEGdhIw+Y
bElpTb/bCbuxxxNqRoD3Uq4n/uEQNSCUxvAVXIYRbZM2bnowIqdF3j7urJHJ4VE+3TST5K/l6/Oi
vO738O1vDNfh3CN1fMOaYJUMIp/q2zgk4t8XiIJ9zgoj5m/agfhiVWKmdM5g4stouW8P/9gc8z4v
jWk2DI2Uh9mido5zTwvrkFtXPHVmYDMbti4UlYgJognJXwW+HCGJqLfcNs9cyYCZ7rQt2JWjVo1s
7BsbkBQCBdjgjq7ZAlk0DCjbDr9u7wy5VVzjywNlBvSltrowq8C1H9jSG55RRgV65DzrtJ2Meugv
JTTW9NB+7ObRedyUlTp2+Xmcuhwma9GzXpyKIaBk8QS9zE9WTE1qgExSBykn+pDQACo7z1GTHVcm
uux4MAp0pFLbax2bkl5gHJ7YVv+RbvNQvqpqTLPNxPRHnPyu15WwawTspPKa2/Z2Rytv6L0gsbz6
BzuXKTUUTZ/wCQmwx/xpIWlAGwr0iiaZYAYEbWI58kxdISG1OJAmQoZaLw9rutsXuIZAE7N2J0q0
chRhZ6+5g2hJW94PO8u3exhn9rT1ToqHvZwATtS0qH0Z9rvp8EAf1NOPk7XmnmzU/+piUi7Za2qF
rH5T7PwCpcPdxCliBGz/CJKYbwIkXCuI2VimwmNjMhQ2jOlY9q5VSyVu878fnVDGvx0u+gNJAS38
oeB9KSUWV4EEudynjlzEIU5lmEmMpaj7PMtCBLbecErDMHeB77MvtSmfEip0bPWIOYNd9vZzjx92
b801CoviOSIQpREVjoUNU00cdASA6fkrl4W1txGWWno9lOTgVKwNpChJp98YURelVC0UDA1tgZEE
qghvBjtba7Bu4nKYDNJBxwGuJpR38MwICDju5DSmirDWt7SeOixzIltUJ2Q6fKJK55MbR/c7l0jj
9fWMgJZbjfor2BR8qaeTwT38EtLjR5kJek6LJEY8UjHvWp+whSoiDDIplx4QmUJJ7oN/1e5U+21N
F3KZ40fnM5dqp1Hi8G0H+LSQKCV90xWeTIOHyOLQOQv3It5L5WHlAcsCayBCIkIFEOjroOh5YLuB
AhkB6gIdrcN41Hnp+nwIG65jrSel2QRhB8bQjhIufvZcAkdMZJMYNHlXBukRE5Vwqj28IO3E22/g
oGXFx4RhdMmDKXTV7t0HKdLyEjyyUg8pkYdUHiCMOz/BrvTX8MwQSinSEPIwuk8ThnTLpFO6uIex
rDAdySXZqSoeXGDuS4jMMAJ/81/2VJEDwKYbmDcfPQPL5lGnA++jrOktkuvFjYgRJPSVJmOwwDKH
43AdRitHJAcFwLJXpNo7ikNopQm51JOc7EYUyhns6qRrMmM2mkWNJop0miPRjZDhJMrJU4nh9pIE
4RF6T8NLWJhYmX+FAq/6MCv6VvcJtbbTSHWbKpnxaWbsbK37I4XO0tE5+aVo4XnHDHy2hrSiOqYH
a7m01VsZqK0Ez58Gppz1cET6rgYcibp7SP01AhNFUweGnH2+m9i/4A/L5o6wNQoOx8DsjBeTraMB
1OEVnzrw7bXJpG91JI9CkVMfihw2BFqd6KDv0KsGl7Q3LuuQBSMeZ5NMiFCeFX0eO98AVyjrM/rX
5fmp8XZUlc4z54fsJzNV6emUBuQ840so/6diTxsHWdwFpXl6e4frCerIW+b0gtTfhAu0oIve4qus
cOolxgH3E/ez9LhUIdR+kgG3/cfsjh/e+POz9USr3sN3vP8kB8jX8RF3bgPQkIaY76P08vhCMico
J37iFnLPe3qIKVJ2vuuYugu5C3urUudumvArM8tFVRuTruxIK/0cJ6Ss31rg/kimPvG/rF+UWHct
e4eI/tI0TTDC1QYWgsHLW1PJES0oO/h92XECYgI1cSircqQuOmzC/NHfCn7svmvHAUyd4na7BDmt
aMZgO3tpkbiQFXbAvCF9NsKFsrTUF33CstqpSoffXRgX3eUQaKIOEdzlMOjRr0YtHZ8QWAAndN0Y
pxqLkQSf5yHDEUpz9O+hnoAD/Pe34B9+feAziBRiVqWUpxGMCIG1JiYg01mNSE7RlKq/yTRTOHgu
1z8yAbCEi7og58L1IkAwqWbpVleA2c6m5QXxWW5HGTxmHDJ0njSeMe5GdVSFB5y/NdYdithkLUQn
QzAt/48f5A49r+S2bKwOhPrcUGAee+HODPSY8rxMcaUHqkoJHmNH+JN7O1LDjTl4+m3rz2q4JZCD
yrjUkvm+4E1l1JMtcrgUai+ufjmUa2mVRjW5B87TBw9curVhMGgJ5PZ46U8vcQKO1I1KI/rizjrJ
7EJxpMwCC6b9lXP8Rn+B9SgCZ0nbGfqKLhVAFRaGjKKf7kuWuDIoszMIVCVP5IKmHUD1OEat06WV
B+4soyJM8H0WA7AXdUYja+XN/+w0aL2qUJ0U0DwTIduFH5xocP3UUNaINg1qjJ10cI4sqpL75515
DUdn+5V4lFcibF0YlsDgdtNXKfUtG9FRKCSpAtvVARki2nb4be4T+QSP39idjg1cNNOVdnd0KU28
f8+mQ4t/NR06l3tg3t+WDn8CYJ8kJHKYx+OOULfBwSiJmHXc0d3b2aJ5Nuj4r39PLScSzVJWbevN
Rh3aZvzYNJBH4TKn9/oYv9eYtZQ0nkxsBHU9j0Ope8/rGHAX/Xvkb6tvagXnJu1FOOFtVhETl4Sv
X8yYOGHIgAP+iL5L1XbjyMpcMvneSYARJn/Rtd3SptmL3a0GYC9G4QRaG4rDpLqtz1WRrjfj6/qm
zrJIB9FwpCsSx3Y75lrWx+nfrZhmCNq3yHJkwO7z4Rmz9xwE0a7/R4SZ3CJh2l94+MWgQc8YUsTS
sKrIJqc0ar/pTMt6bBtyrxYw0HXox1RbW9cmYXp+947gGdLYBTo3EWGzkJdbaj1ijR9pAgYsHDg7
wsD4eOeCIJVBcQPVUMJsyO7U8JbwpJiyaxPcVPtGDvznk+vvH1S/2G++Qu9oeor2raNlDYBoTN0a
L3onxvti+vxMzWyrPMg5THjtx+cH+1jE1tLiMHepFRTxsne2IgQVKHPpQX6oRx6B5p2OJXzSpYde
d7i1wTLLYbhVs5anMXRicbMwckdRw7OdL7kiBZFt5cKJUAG2KlO2O+hBgbTVmuV7B/Pv//ylf/F0
rWD5TxF/8F4pPkFDlpzbxiAjesElp8xUFFYknQ/tMgCwyeGtlzIB5qU/8ygT943RZktwwPTJMAko
Hl4j+gWrG4orRzx/8Ifm7iBaHgJfdncYEIiQOm7ck8jr0xxRYaE2fNAQtsKX54R7yySgCH5GRBj+
fh+PCQZfz2iP4Xjr822OJsFIxs3zVW13k9OsoLNwWxCij1eIsWnzFIANUfYF9wp9q5HUDmTpT0Jk
4pmoNatLFoepjSWY2mv63o8TMn3+BeckmzhuubZSEfP0un8IOviD2Ho7MdRt92IXt62s+VitRZaH
bWiMcks9wMiBlNbZY/KNL9PfaUOFbo2GYpqo5NojVNn/ONT/oM3FRCwymXS61FrhCltnFghuiI6h
cOToQkxyqgLv8zXYLeGFV9hQ+k+rhNjXApwNmMBey1nJX/F5X9qir4y/twiZWn5hMsn5Goi7+78B
hKdC0Q0mprHkmq9LSpyXTDcE5fOXwPPzV8HPlahwW8RTk1Uw9xderNrSoBdfdz8zutDn7Iq6K6j4
bLYVUWJ246yzOWaJXsRuhHQX02uzc+pQgUlWHgXrxDcDyWS7sYOL3MwbGQadgo7S3WQquEq2ILXa
jIEMo+ETjE9EYV2MEmGpxMHkjcSa+WqYDDos75B6JpD+PAdAr00Mikios3/kgN9VeAlidyF/2Xxa
/qLNZcxvyB6SJc9bZNXlZiTW2JL81DRM4jXsoo/HdV4aICf8aysSYito0/qY1GLT3TXEIn3By3GN
QRZnROTxi3Go3XyzSmKg39YcCSH+Ktv3lvoXBXEECUA96C6yC+KXZOOzIf/iR0B+j0SwDnbfFpFY
TJtiF4g3TI2s1aSMVSsrI9MQg7Yd4H5+r0Dn2a2QElWdhjXIfwNqUN4lLAXiIgCa1rK5tte6Zdld
uCIuNZhZxS5AB6eAJItwSyA1DdtiS/hz0/K8PPDUKISxTiJf27sZY8Ew0RqjGCPYyn7FpxsmEOjk
YV6BlgG7TXHQ+vnH7Wu8MVbMdU9faSCSTsqR9ELthARe5BT2WvhwEu8Sjh+/98xhou36hgnfdcTb
Ml+2qIqp7+nKKdIgH5FiB9PyfS2JloqcJhqheHb2v1R1B1dSemfeA2PAw2uP6fRviS4eZRYoW3f2
cSCBCuuo6v9zEtVVdgTbUoS37Jty8LmDjXJQJfgySqWpW3wl7W5djfl4X7VI4gU4UY/KtRANSUCj
J+n9tUueZNwd7eRngNQHzE+Cfh4zdlOI62afxwN0gmrQBWMtFxdYwgy8GNNJJ012qQBuujHP/ST9
NJkD8X9X/4oNMNa2ueJDW2DYWVkgqjZCqxH9rE2LSJwiI1MqyCPGkUTtvgF/yyyMROtesQDBkjWl
y/W1dF/Vx9iijg/6+VlxUxAH6335/McNyvL6gBOVVPwnUdYeu7nvu4cnLKP8+B9AwcCb0vz/bGTS
Hl1SwpaRx+NS1q2S73XypA+8tPVhZomrlky4V72/UkEAcd7QSgaAAuSd7N7Q6JbhX2gp4luMGj2o
B93dGs48wJ5nIvwq9uCpLtWxMHbNUshvI0TKVD/GD7uG0CSJ650AvoivJ401oQpphewt7lgrCWK7
1d5/P9BUM45W5raYLoIC5VN///FKfHtmeWIx8ZI756e1G51FjIS1WuKgoKBIvTAyJJO8OKt7H0K1
tBn5VmlK77Oqs1ogCYD5JEiR1FRJvYru9N3BpuZIrxGDJ1OislKWtUqW5v3u+yUI82pzK8tm09kv
y/nMdgysZ0d1njbhK35tJEq6nC5RZN8PmPZZQQL3QrRRJzQAs2z4wt1pgr1WgHWHlOwseVvLU9/g
a1NJ3XteU7QJ8y/9z/ivj2uAAHj7iKAZ+hBmyRQaU+StdPghxu/0wlYCt5D0K0OBFIvizfpTzcY3
InMNibvZd03swOt3swedJHhwupRytO50hRm6XvqCUEn4JpydXFW0XMA9e9VKVmL7Thv3dlZ2RZe5
2GFsWxe2J6VJO3eTC5QUnuq4ARHqj1GWpoeoOK7CNj848J6EhFULD/Biag5x0/9PjFrSRAG5hVKm
s01UEtZN7IqNAptwrSO3QPzewllxirU8ByMLzY62CntdUP0HxxbIbgsjLqFRgopXi0PrEfhZUhDX
lrYWLyjPlZGscMtyDJ9F6JZ7BU/fvISi3EueZGi2NbnFHcQMPqFfIdkvEKNZMqnt8Nfp95yWV9nf
tuoO6XInPfMJUn4f+i14elo+qGjLAnalL1cZfctAkkn6e0cr6YQNImJBGHuk6s3LpcJDowRecJRO
Fd2z6OMflhTvCyE+64rpwet199ihD76kYLpZkwPnxZNmegoHhnUx6Yzna//SJ4m33xHIZgPR//0r
FeBCeJsnfHqcEx/apT7ua29GgDsTkG4oKi+K+404jxfew6ExKdeamHx+19sAMjPr4CtcjaewR/Gn
Qd70RcLeZ0UcTGFAdieN1pLxESQrQ2dKoHh2VVgILX1LH5HSNn1YyY77Y+cBR5nDbIARQWMWSYM9
bgwWnDczaDA09TubjAbEHm/wuA0ZCp/KhqAx2Dvduf+ll+PFpjegSTrUTEXx/gWWgyluEzjeucie
tJZrmcgigWwjAA2EWx1Mpb2jXPf+5IVd+/0UjTjyia0ZRQKjRPKR2bRVZL7kcQ9kEWIXjvJ9H/9e
gbQvuJJ7dLpUxwKq3RDWtRz1Eq4wkRHIOy+32i3yLZeZ56fjDOZ/2+8kESaHiBqwQkWkw3NdET3C
HzGDGDb6v9q0vP/g8CmCTL7u2T04xiHWI7f+Qg7wZO4FTOhG71HYq0Jhst3aIDF0ct4rRfLubu5h
hSpkEVJCQruK0o4IGavi7wR7dabpb3NhOmBjmMcxQUnOQpwcGJSUh1saNn8oZTozrer6vamr+Qdi
HqFAEejMH087UnEBNYULCzkMaq02zswtswzvjyCn+i1SI4YTSOKBf02CILWUa9zL1Wuuws6r+p+S
eWBYCDXib43+UBzH6TfHmPGrS9w+V8Rc5MPztTS4JnMJpNlx+uwk2kEPeEc9VIMJsbh3pYrNEMR1
KHI65nze81FDj1GaX01bVA1aaE4aTVeKIzd3iuhgUSfkUt8/npn2J6D5ljYiO64m6g1UrFh2Odpf
aMI/je3n4xvA+D+dAEHpfa2f7MzR0+DPKKJKEYR+KXG0g8IO7AMOOtV0EBVRVRopS5rKvts3RdMh
4B5RVJ069Yy38288gvMRNWhKMdTU4dkFvlvB5rjG0hqmHWFmj2wozLzcnrYTiwB5It6s4WEAYye7
V6A8YikovNbkLhKPtSrruQ/EFjiC2XXskYAdyfSa2t5D0/IjzeFhJhc3QDIvgkG3YWD6nA30Q0jR
Q6KOX2OJA7XO78gzctw/ZYtHWSl18iVF0MkNvTqhU/oSv6VpGfQbqZeWYs/n/LQxGHGk6H3sugmw
JMenNrlblfzRoPcxUjQrXdjsLl1ohkMeLAX3DSMMb7PJ4Z2BB3EOuSn6rRuFHudUIx6iwg4vKLAo
mFNlbMOgLVuWfnNyNLYiQR/S3iX9iX4IPRsDk1XNf61QRaQnmy71dfIt4AI+gjHWaQerLUTpgeWt
1AgUxUpjp+aF6zgeMDaVS4SUBuSTgNFiJfsqYGAy/s9RSnqtl8hh2SMbEYB1BRa0Sf8RUvamMcxR
KNSO24VAxS7dwgxUFGvbjaGkrxJlme7RVUCQps7nKS93HTXiBg/l1n3rI1RL0AWYTP+Dx5wqOhzu
OCBp6TD1hWdK3h8zPzuKz46adAShtJdkwcnhxcHhha7rBvFkigZhEmbQaS9D7tIOMGHbzgc3Igel
bLFiVFPAODjMANkNohoG54BR5VoGdGJKgCpEtdobWNar0OTaE0eyqe7Mxmb2bGM2bSn8beY0Y1qY
04WLWJVNbHI31ycWiiULiVEysIe2Qemr9Ov7aoSl48ydzBQs+XKC5t5eHAzbcf06C0WYke8SCJTz
mw5CkyRGrak+WlU9oSQ2399MotRmeCqHA0veGKg7MI7vg9YDizh89NiOeGOQ6nUQ1l9DNGWfKtnC
cVyLHrXusst505IPt/5K777QKaQGv93b1Ba1StShkS2dMYAJf+SOcA/RiNAj7RJrd4jL6WJ5DoKf
CMtNrGqHbCOa+TXR+Ke6Vsj7rvhDMYvfNP4+hqSdQRl9B3NK4BSCC6/0S407BFhlILRvl8mOuFiy
vSNpkCG+9PZxXgYvV5nvjHkIlOg4oFrafVYDziKpkXrDP6D520wmelasWfAk6wIfqu/GlERQZ3N3
/bNAeoBT1V83P1WIR9+058tKwrcLUQS0wuqxC+N9gcVnP4MMN13s3esRy71TzNbkMzhQNtr5IB99
QPJBTxnve034dNV8Qn9tx/iziTyGrwH8AkJW0GqZUCECviLjc0r0PPcIuUcDDf/Z+J2+FNdSLVnr
EDL60XuIE1H14vUT43An9rltU0i1rTO3t4XXpyTCWPip3MFI3hFSR2ebF4lXxtmS0+F7PN8w2CAO
90rmEbBB5zjahd4gqyE5VBTGHRUPmWWVMihyQ8KpAkg6AmWA3wj8nXfFAZKEF+CkUcZu7jWE6KC+
Vq1nXzaD9PrUGQMVVbQHN8iA8bUR6zvtKb3iVOzisQGDVBi5yNSud1L4a4zTtiuPijYs44xLR8Ik
1J31bbziLDE/M19YcstbtLNkV/8Cx58ZwXVcUcasxBHCGHb7tnySROz4WVn+z+c3Eyv3LFE+QbKH
kfoewhkmeTtQMdlaBJ/ZYgoMXPGEFoq3x9rgIMRar1jI9FbFkLrjiV+kXqHabkrzrIkmhaqC4FoA
4hJ22YP0PoDi0QhmY3hLTamYhUXvR3KfQMNtGiKAjyJAfK31Tfl/3lJzyOTzZy0mGyCwgDHp16AY
YY7ihgk74yK7Gg44sj9LRXDnC8ZAuendSWHLbnCzZY1BnmF+pIGAQ8HjcPYWw7A+dRg0ictr/fDQ
UVzP0f9XZoLrTUZHn/XwYgVwzUilRy2awl/ExyqTOSalyMh77TiwPO1z59w/3mt0RkZtno5uGi3h
DmuyenRGIEyy1N6fOYLrezYaCeH+ziMT9T5nt+BirFhNWVZTB0DC+xXsGBUaQkdHvhb8igkzYuTz
Apktu9mAaaTqSWDXdmVchBswcehiXh0S0guT7BF/1cgZfyT6c6mjsgQVzljMU8j59hqLfzoc1pc0
2flFJj+igAZw/MDEHtDck+tvfVyz/OHZXYiYjXYMp/njE59/Hi2Y9E3Il13e/5MasZJH26wOnp0K
2eluxcgDSNoGvbKehNDOW6sJPvnGZB+JGG/wo0ZlQHK0UIi8Vp9BFrGBxiLf51vfNjyP2ZtrltFA
YlRGRXwuTUp0QBVncUoZBzszFcDuQt1tntX5loHCfD8NKw7XY9FQRBI5smJYjGFtUF39VhPDHzAt
CkEQKVDGCZvOFsZTwdwoHtSR2/ErlgqN01wYMgdfTmL/zBW/n2kFzIGSJrW3t6+MeWBRBbRQArQk
FVRyu22bDEq4+KdO9qGXw+rKMNnYx8jAkIuaTGWANbvt5oTwCDegt4Z0Iz2TW8pSfojaWmO3GOEy
sMYzmGZIzJ0aWEtz40ABF7lbvbHp+xVBX4SpcBdwvLmr1zBHVKhK1mrW9e3lmdF3I1x6vqEFh39m
sf2X9WqTUhMQfLtA/2vEBwi5by5+addTSKUYSsogaxtNao0QYT1wRnR/MfsmImDDJJRohG28vypK
oWO1r6C8qd1fV3ZNn/7IaAHbcETijDsJidJHCWjNkZrm4uTHFYx85GH7yN0wFkc+nUe9RkTG7hAU
Ls1s9BKquQiSGctwee2drxJ+gwQG/V7nlZ0hIYMHQ7lfVU7mmYzozUEKgqqzi8VT5YjvCM82lbC8
g3TRpXO3aIbS3vXdAbjcZgraiwlBhwWwMAj5S8ngCLz1rOSq0vqitfouSUdDixRlIWmwCDmzrTs7
LtT+9hNdFN66ZeCnIwn23feklPXfTJqeYRSgM/yp+s4VkAa99MjC65iwI41uPOUcm5XmZzQfN+49
5Vc1uDWug7laoYD956+mbof3+I/tzVcCqOjT4ugoqK1cDTiwORVJR4u9/7sDBGtAYkYNwXciqD36
BKiqxAPg7kL1btFGg9Vc9sX8fzxiI+WcoZnpPF4GxhP7vGHJD8dS/LB/1OKSR1tg0qyuraFdtYk0
LUmN0jr356J5VeCQTs5V+EMAii6x0+d5WM4cYTq+csBTJGUbhMzo8PiMT54/T1Fb3RzkfdIp30zj
QYuZOuRZ1lr1fYhQCW6QReXemAkWdGDyP4YL8MMxkL9PrukHL+s/Q7O2nLuqWImj7T/PjwKupBNw
wJlTs1X9i6mCqYAw88EcSHXMcZWGeOmsuyVFiQvF4qgzCa0D7D13Bs2ram1FlrBmWIKBFy4sDZSZ
YAgCkiZ+vFqad1pnz02Af5A08IhxZLGvOHLHix8JL3hblRmULVcdAYHphCxapr7Jbwmymro5ot9P
rpqMnbZD+RXr+W8ik3T9mtB7iGUJXa3eHutfnOxzxAxYbtiIWoaN4P+tY87c3IZhm03DZ/j3GIQ4
ohkH7CppaqWl4gU458m3P1iBx/JnUHqlNQx61Rr+MpEhLlNkjhvfvlYtCuw6yXfOmcWAMs937vqS
5FdjT90xqYqv8FhlqsDo/lfPj2J5X6/mAG2yFYVwd+/J94D8qBu0s2TShdr+rDec+3E/Orom9ktW
5PcLgj8M0eZB6zC8DqXg3zqB50ceGt1dQ0r8Hfet+nsl9OZkx8rZbecw957gGiM8kwHJ1zudJmpq
VW5ai3CnrmDZ3LXmQr2vOaisUvFOXMLppCJ/cQ3MXbGe8jedM7uOBJZx8zXbGFseDy0J6itSfr9j
6MXK9967BeC+6EVs01uszFE/FZcOVqRQ48DdQ3crdFa/bl4geo7JXT+z3x/UnZruqG+ocsUnheF8
xjD2vHNANkPTY6YtBjBCdQSZ2ErSBTee0jVmHTOVZR7l1Ha5aoAYWLeNbttNCBt53A5vERQTb8ax
MeY0Kfaee1/AqV/1dR7oIuCMaqNkRfz1i9ponp+/sLwi5SJtqHH3Pz1jF8IntF4XRyQRUOy2m8P3
ZYg+e3nnwW3obTYZ+M0UnFeL9bMU3ylPAXJrg+ZlqcwynXE2kTlVJ7KAuf9zvGbV70CpYIBS/t6P
Ooa20kuEjh5oFewkIfU+zWo8gTk0zQeKK/Tt8ZjBjYqqh05HIiFM7IOau4+ZBRmEmyf/fZvbgimX
yAuAwoqwJRGktVI+VBObS5OITuu716O7rB4L+7BGoBNmD7ILFK6A3Ksf+JWFw/PpO0ocLHY8H8gN
HOrH6ZUGGVN8DpG4aTRKTlgPWEU8e7kCEQWQGyYme3gLV+FbI1xS97vHe+iBLDzTOFC80NG+dE1t
xLNj2TGSMYyy2O8sOaQ+tMkSc1UqPB68NMk9DGSCE7DCUSd0AAxeK7Osmj27xI6JhCnfuYmiD9LC
WK1yoXtehMwu909+/3iyihK0pb5BxQPG2eN8HJnOl9uw/bjEOmHaVSTo1IbxV1cppucg0AZW/d9e
ORYyV5mgyMfqggMdte6gVixhYvqOgQXdcIwNf6ml9krm1myO4O7Nyr1iB/2e2crwuthPQnTMV/Du
853WjAZVQJ9VON5dLHk6h/auWAf08L3llui5K6JF25zbXzSLq+jo/+XaMQCM6+eDPLeeGb6xUINX
w6MlBK1uYXfEaUIu6kFhlyzuBPgHjPUj+aPAZ11Jcpw3zwlMGava2f9oq8BUV41LlmqcRzbZu/UJ
XYKCxDzpiVDIljZ/21Vj2/Sah24Kce8sUNuM8NbeIspHTcchkuz3G84jCYm762jIcZhgmmShwynP
IkHaD/AnylI6Fz/x8yJc/SmGLwyI3OK99fG1olvKAFReHLeNiJZ3Xjat/po3zfuE03WQUYWbnq9F
tC6KvpxCfOuPk97nhgAwHjcHhvJ3LyfZlsnwlL6jUs8amQ1hksI+Gdsxod1amoG0ZQZygpGzS1cn
Wrnyo73Mjpfdsm90brv8VzP8frIIJLgiihnSq5q5govdvxCs0GWu97uYe5owi20aZk8a+Gl7Q6hK
HoPI4eJy1K6/D8PCimmwrmWGWH4O+8SozjYb6ajNM1SzxvEv9NMRicjte9VcKgencdotc6OXHF7F
u8qwF7FZB2TmU+yopLWkJE1hnRQWkjZyGJSdcO1h9RUsQar05yeDyvZ3Pzws/aK/t1DNnsDZNt/D
0AiE/XvlS8B0w8i/UJOeK54VFpzxdhclL6rJ67cWe4kGr9uULfjP4z7gp0wW6o+5DlFH/HGAHdvW
+IkrTZiL0BYFYpcpydhyJOmvaYfj9oezNh9spc+CsG17x99cClcgLUAYSEn83Vz5ACbXrOqYS0K0
tqzaN+/LudjaW8TywBsQcOz4pE/nF4PWvNzhY+xYD11Ip70vrQwhgyIW3Z8dQ9fBgZxl9NkxacmV
oWdmmHXVcfVSq2u51FAM1E07CWIuVQOozDfucaFcbIVFy7AB4ZnQMf3cDBMhSkheck8jXC+0ijus
3/hzg0s1BWQw1DXI9+Kkob5IRMeIDlneebgmiBd5S6rD7b3N9EYC4GFAltRpU6koYDFPGKPiXzNm
z7VsIHEnbTYfxqCE23koJIj6qtDkF4GlhaBmrPSsyNwBw4dFHs119LTamu1ZuVZ7O9VKgUxi2+JZ
GwmPXKEocEve9+Hw+QDl7IIuTKhOmWGTv9pT25uDYrXSMxBVDrpDB/odsJrC7oexw4Pw+OnkiY/j
d05loeKL5sK2dZUA6R0n1asYXLp3hyKi4QdmCFHJbf0T3zSOnsseyTbNQfE5IniiO2xM4REdIQXE
RjUJZsIxuqkH7V0yPG154kDOMfooCTBo7oqODicNVACoT3Deal60cPnh9ta0D8RjDtelTcxK4PKf
3myXmjptvpztBsd4DH6HCXkXuoAV6lwkrdaPmPW+1PdAmPJfT25X76SLv7yWduWUJcozCnHyugd4
m2gqVGYs0w0xOWM9th6iTZOmHMxE17bvk8LcyQCcZF+4WDfhf8aKsxPqcus5MCU4RBqdEY2J8619
BqILGd2FHpv8O1FwWJi6zUhskLeAVmY4Ga9i+lPEbEvOIpiUxJQV4aJdhdT3HaW8o9JaGYLx7riN
l8rqTRLuWIX0oRj2e2F5S5FWgQSv6PH3GNm3Jy69nTu9rZefZ1/ynoycXucGvYbXKStvjwnJJPhd
PddPaQaZPUvuqXTFvhrX7r4edAoFR+cbORUz6WCpWM8sLAp8+59Dse2bJ3heFqjzA+OC61YB8oPx
MUOhhscH7pzGO+oBMAvJfDDoFmINPk4y8vccQouIHN1bc1OSW6jljSQGPDuZn7cqB96e9zwOZIJm
MtNE4f+Ga29Uh/RCFedglPENAZerETfrvTEtyvmQXJ/nsdMEiD0Df9VKsI9/owWeIElgN5hdubdt
YZqC8rlaoMBTPsQzbJfvvUMMbyrvjZmPP/0OwZBEuPm+sWh42dT238ekgsw+8ZM8b7jSgb/3gUGH
jIHjBgfiPjBfScOjtylgyHkUVzfLrXf8KPoGI1nfDK8JesQnY988D3tMB/8tOI+rvPGM90aJ3bEM
71XWZy3AxhEuNQF0sLBGIqJCt4JnPHcEbGkxHJtUwjORvsoThnbbXUoyIIzbx11nZu8IUcaoyDgm
wSAhd+O/COxvCdjc2qkCTilZIWagukX+PJFFI34MsmI4iuS3kpIaSITtXX/0FK/paLVCrc3bsgyf
Y17RZQ+TbXw+x3Hj8pqCuiPP4FyzQi8xpXVZcpVb41HETxmbvlKJrkqxsRt1/Isxswz0w7Z9V/mF
NpgzE21vYBbCe64VIkO5iSaHIqxLIeOZpGaDzWpkBmyGxM3xf+FsGyN1WckN05EuI3Upq0ZNL43r
hKK0G2ouxCnOifwE1vNp6w99Zxi6NNynhLrAvupc9RDcc7th2+Axu53FaiU0DuEJ6an1pcjOObBs
aEsUT3c3fwKCBtPos51YySQAUXN/fCL5bcuLkBpe4buDFFSL5m+rwYTt37+eudAZKqz6JT9fbw7n
EvXU/0pmOS3scaBa3kdOfDX+LJq3ka63xfvJT9uX2HLbYh1vmNUVYIjr544snolPtlJdK4X3bnpY
Ic0gjBX61i/EX4JPu1De0gx4ZMaxhjH7hg9EbDy2rDbryJi3szn5xsUSpsK5RZJJJfjBBRvjeVwB
xD1ULyduYoCPrEXK/AlTfQ7d9YH4yjdhTULmRHdzE30lVcrQgazNWzZ6vmWx0Sk2xAYOT32rP5kV
VQbZXcUxFcjhmcWqq1j/8iTCCzWX7QiJp9uzVbxsV0N/v3dMtnOGVI70HcnDJbeSzThTPbK8Cd6M
KindaHbwU5B+zpPnUf554RjfNeLb+Li1cH1nE8BCKBa57FYcp5jE7IolKtAKr7r1bNHhhqPuVsre
k4WRbEG7Hg/0GFlgWvjWS6VCz6x7NoFM7JRWcQkVo2MpjKybkNhO694Bc4B0QwezpMoGAY3USBdC
AGqeL0MJO0djHfb610Ed+2I/VmdHMQJFwbDqZTrTRZtq0hsTvwaG8lV6jMzq8D8G2nw6EnerEWZu
eC7KEWLeuu3dy3wEMiftlJrWu+FlSgTSIky76/BB0h/jvKE87CaFTFabri55FFvRM7wQ/0fS8Xrv
UMvERJvdy31B3xTDSlX43iTQq8bUEK8thqRC8Jwy1VaqA/8Ym4n9b/rDAGW3ExHq3S3f/rHTqN8W
Ub/Kvym8Q72XIqZG9jUIw7M/ihXFl4d3biGLoMzGPRu3ZxwlAIXUdK3A5FYdfsAunKgMRzmLBxQ+
cK5lZMNmpOE+JtGfp4ZtGQhpS5UECCFoK4UDYFRgPO2CEwR/1qLJ56Fw88+o9JeZfMHSsR4c+1oD
//ytBZSfoLVJzplyUXmBQbQx+iRDXPIktzpsnAItb04NRWIBmZSX+vzAFBX3BToJDv6ymwJ5Uuqe
LaswEB6gDDgt1J+H7eIbxZa9vJN2dSc/pcJwIh61k64uT3bvb/l+C9DhAyQ1NqTTqCV+rXv1Qgij
WJF+dmT9g/YFnHxkIbgpT86qylViFtsLulXa6eI20PFZa2I/xNsJC7M5ITnA+imUpU2TXukx8ZA4
n419I+37Furr0MzcFZB5wq3r+I1AQWCX8XYepBfGo+8FVHz8SWj4zy9xynICrz5JG7yWFaYuRhl0
vUrX+N1kRhmaQqI96ueiyA0yUSDVyPuM+7nyruKXcjaxbjJFFO+5VjQFJBZyAHuqc+SRmb7FbByw
S7NOcc+KLmoXHgffLofwOhpYn+bnlcB0R3AcJR1+Dh88as2/Cy7seUYwjBnTecB/FyRzhzW5I0Zd
HLFizDE5/M5GGPHEYw+kGCSbqs1JcKZyiE3iAU86F6lFaSvn+dz8Houa7xqCOycN9QY5QZkFfcsp
Fh+dfvQsqszvM3O7fPrBHys/m4eiEbbkGZMRJvWVUaMuI1m+6sBApDCX3UvFS8HCr3kxVniCVe4m
KialZzDWXxmHGxAuO4tS34xwdIo4MvVl9mEakOfepbddcBDG3VXfz/Gwp+IGgOlvroQQNLMNZIr9
D/vPNQwiLDtsTO58DllyjMM6qzgYmQsMY/PTVGISzShMC0d7crgC71vGkaI1PMJuu2Ocg60zS18a
fwAiFELYjiMixKXd0aMDN+jZXbybsA8f7MkRmT48AdAk3TOj3ayW8m3H4GzOD4w85WuhLw2rA5Hn
2XHB0Ffm5KjfKv66hy/HZOT58sudFi/eNWAQa/OEnsnrBsx5cRanr4zw6fyphrqcJVQuHOGj7IJt
gchQCrLlrILwIKvKXx+c//OJFfkwiJv1+HwQr+gYDEwdvqHNklgbFysW9YSyrYAzjuCMfc44O8qf
gjZgiex2mUy3FWqQWoK7Pzemh/kgSl6JgR02U9iQ1jScje9VZA/T42Sg2sRC5k564VxOV7RhNClu
4BGd5lzpl9aspjmu6alVel4+CUEJ9Mrx/VMtM4yRwqQaR0/GuhSZUnDcAlbVR5rR5G6tVC2gtDzk
eMURGnJeD+PJ85EBV3No0eqRLf1nCHxraXbydhh1RJK3vSUIR4TRVn1jKMM9VRhqr/iI1XEmtl55
q06GgCABp5RGvuwp3jmULPNtrL5qNmZ0LcurLg4zFLpCrvx3L/6hDjb7poelh/kWnOyqxJw98g6x
XMNIP1S8xFpJXfMxTDbdNeOR6xE77Z8vZXrs3Obfd1W1fp2+w9o9sTVAQbVEaMPP/Of9ZPIKncsA
oUs62zoppc/Gw7dZsVOQrGxVK09DjN4GM1s7ZGTpqsxm5l8GeJ9iG6CeNlJtfGgj+T8Pnd2hrj9i
XvL5QR6/sIQ4Ld55BGDd8AaB+XMuC3be1RPYpWG8KTS/rAsTYWXgvJKwbkDRzkiez9ItUXRctSu3
EqIhz/A8HobotHKbrZR6FRDaHiDu8bHFostgPa++iy3c4UlnAhxE1LyVqyGvrBmuURua7KXU9KJX
3Z1VooBw0lEY0pN+M32KygmKOHDLPS5Qv4cwpYIqC7Zho+3K7FPEKKdyuIWjMLxYvV52+/eY8NOu
A6/6t06D80/EsdFWu/v0WSOnyCGDctdLYT+34penAaRrXyCWzcDkQn7I6rGsvfJii/tV8eDoEZaa
IZJHCZlsBGAnE8bsaRIU/YWtKOls3pcAI6Te5aljXYHDeT3voyWh1Hni9ZvAHJZd5c1ANYAAhO7F
T1g02aLa3fx7ak5sRThwv3RnSCRvLwpkEYoKb31Cnt2hyGIWaDAMPDkcgMPyxMpjfWgVQbqQ/8wa
baFcBOKUsMwz+X+mmM0BOeT/aGo+u5L99B8huXSZ7g6wIrS0mkU1K30AMaw755YIIN72s0BgiZ6i
mVl3s5dfr48YjOkUPbstfd22Um/W64Wu9y2/tLT6M6qAVEZq8kKjS/oEYhs6tGqkPzP9ENoGMsmh
+RdhgPP7AYYItHqTovRt5RAdx5XVH1Pm+CPPqta4gVMJF2xfeolElNRi0hKH/RhMKVmU0s/bbmUH
hJt0lVN+SC5e/mbjKqy5qYp7cBU7JC36ajad1U5ZAiexoalv0TNIfpLL39a3kBfaZ3YyelnyoWYb
zEfPyy/Kr8mIjYeFYA0fFYlL3Qgh6aDft7xXZ7fyzz+K1mMsdL9pyXgG6yLW5VCi8vrVB67PnJgh
8rM5IDlWczsF0tpcouB0ZE/Cq3dch9vU57nEmyEnImee8TPcBm9KMVehvxpqziORzXVBGbgN7Z8X
uW1GPzZsNDs1ci9lmK/aIsy2VcH0Iv9DDaWx92Vnod7px2uptni5UI/5M0EDjizyJnAxRhE2a+yt
Je1wle+bwXSiNVxzirkmeVzN3EytgAGBlqDWju8Otn1Tqq2KzBVwHV9NndHprJDcMuUSV3lAFvhB
5QQEj4YYRApjJLy+Dxw38pwreWEYs3mUTIB8N08GoZ1NCINz2mpFxDkcpb5G9RHLl3t+6FhvPiOx
DDmpOjdmv22EjcJxjb+qdgRbnc7xxGZWCBEIPmPHhXx6Id3r9t6ipuODsqXHLDzfofz/dsaE3GE8
Cm7MgvjWC2eotGfzSdpT/e/vINjxq4ladxqXgASnPUB96RaS8aqWWnX/oBJkWJuWm3q/rT2wpc4G
E2UbYp8hcKe+L4oJyLpoWqzGMZyToeEupqIgcHiTKXlJ5NCPtsMImcrim2AQ4Nv0+M/NaXbFgN5W
oM0rDLpcwevHRnZsvMAe1QvDAkZaOeS4YLno/sTDDSvBaTsFLDZfF1bJ/ld3HqU6mHsy+b7/NouD
7YXELgkvVYP+lkwwMJMQMiumJBvTAEWQ3SclKLK9TG5Q9llqXeadXHk3UdGYYJeZ8dO5haxUJvPw
oVAGhnQ8nccGLM7FLVmDGs+QqKX5BCHKLa1WyL1CsSb3Uvj7j2fLIY2fq5s+jpWx/R/8qJy2VJaG
UT/ky53BmsT+4TP9+sjAUivQci1ck10KqTFEfCmvYr4he+gdnPAPf83OyfC44Qa2FeTmNHaEN4lK
jb3aO+GP6pm9LVXab8uqN/Ho5qgvcVCABfyJZKFWVHoqpA62nIVkDGEnQtHlsROqXO4Sa5nGX1Ml
qdIzX3RByEG1tICWUo3kCYf5pJ0+WXPRR2wUaPtMc7MFeOPAiJEp2xiCNmq5Qpzosg/eyNCe6V+j
GfxnMCJ+HtmyIHDpn5UJaOifPRP/V9B5sLn6I0ssI/35sgvs8Wvzg5g9rFRWv9roWL32G38K+tuP
GMmWUoo9MsQMPFg+h9VC9qVGaACe4rqMFG1pRfxUiaMMrevFYM93lCgyGs/YZ0XBY4ehc71Ttlib
fuZkWmnbLbcdqVglfHZAZQhuS3EhhydjQmLU/xulwSGt2+H8h3P0y2e+uIcnxcWXcgmDPlHVZrhK
HjxvGxrbfeoUbloXrN8/7wXPYwarQ/c1HEcUGe+F+qg6iu2C9UbovqKLPAmUkPK15uQhfdTEI4N8
YhxLX2yC64Qi8gcetR2CZT/DfLXNynxVf7rAebxqCiYP6aw2hYc8VwpUZwunS0lT7NvUwhI7XGHA
LpkYruPcao3CVWUK4TxsYtnKp/BrSBxpb0gfUBdzD4AmCg8FU1E9xNNouSxKErVwyFo2cgQBWopk
WRhV8S6udH+VnpqEI1tfoX5mpcn3dq/fMDRtnlrvnpEtT02sC9pw94eTT4V2N678G0pTZVBNNS8k
El30gIy4DVfR9mmMqDCI6PvRBd4YN4nCn0xOUX4wl9N3W2oCH8HffcnfyloEm9jS7+FOXQgvnMHW
Gaie9lBgUevF6D2nVdXa2aeLWmtQZee+qZhx0+uEjUlowfypwY4YF1dsTJme4K8Un5s5/HTvcIe+
vN2Lt/bKo61K+dm94Jodm+GO3t4gxSHw5jCAsapS0UmKBCeW0TJymqe9ru/MvWvYVnBwMyn6Dijx
o8Gh54ycYtXsMB/NnE2wpEik0jOlIBYAnj1eEugUcN0AH4QhXPOQqYnt+Reyj4xhTUE/9CSPldmo
ocxiLdLdVscrz9fhUROx4p/GZoCVvSg6XbSMa+WMx9FxWx3huDiUp2jerZNM5B3op66fCiwRvmH7
8SUVpIvjTVTV/m5elCNOVlrZVjFLObHE00am1xmY21ofpaufFTpV06lmJxtdRN4EIlYjuXO8cUkL
ah7gzGet/gSfHRZQsE5gZJ6V6yUMWzP4J+c4aHl1IJuc+jEiNDD1NW3tFr0wiT9YBHBctNCCmtAQ
aMW+M0U2hW89UITDW8/SrqPPzeRhEpGQJsxv+v9Q87gT4Mcv2GuUfp1jiEUXvKB2m9EAIwxVdD84
fkzl0hOwDkvvd5V3z5nC0us5rDSVKeI4KxrUq4EfteVWU5nz4y6zYpb44QjsJinNBQGj6PCY41uB
2cTaKjg1bOVchAJxFsdzzDMjNsUmFzpoZr1tBUsCBFevqjbcK0d5oEHAAX7Uxf2kWNbeWhJ80tzv
rB93H3FhC6zbW72tjsWZpCuU73SoMUozXsUvqeNyGZ5PZhWpTZY2tpFTVrYpDNfrGMHFk3jTzw2t
H4zc3fQq5g15tvNdGUlcArDBcctmw5OLONY6DdJHZVkADQnX4feGv5ij+1pqS9vHVZNy81mi98SU
gEsUc9eJkQxozKHvA2BfgRrdDvmRG5GZAZT7mQFdTTCaauabAxCqSU9PxBBb9P1GuQJxG3l256jG
LM/o22PLgt8VZ5j9cksuytaD8yKxg6XU0RB9nh1CJYv5Evka47ReU+SYbTeQOa6X/OD4kEOmMemV
Nb9asuGTEtOeLht9kCsx/fpkwbGA6rrJTwyHCou1SzQDvMxRxjFi1a3dlRUBO3y3dZcqvLyZzHRF
R/91cULGMs9JsIF9P4QO6ED5yAjU2MsamQsgxCnL4a2wSG6+bqy1RUI+yHJ3FKF7aqSvPrFF2CCB
yOdo2S4KORS6MSYRxORiMrrf+9N5xXWX5sNuTKhcsxBatMQhCQYC0W/4IVU4NJqVNXIeSqt4fh43
lwXb9QCgVjdWwZ9ADxes3p59CDX4atv4yPm4YozmzpQQ7Q581GHMjL7ZNVrtUXWtQNuUd2lny6QT
48Ni7cxoR/cjxDdfGWtQoz1CIvPNMczTNV4S17IHvdM5Io53Gq/04k+ph1tD682DnXGdFuGLOKtK
yUxyONWQ9KG4uD7sTK6yIKLon75OCk7qf4ZbCA3dDTE3cc8+XTYLy0cl3BxOPST7zYZDE1CR8I3T
tJsy5O1SMleiMmeXIyM2I7x9bygk4rlytBevYLIOyVYFbdvn2+BiOqOrzWdvSjACJn5a0OXHrQQO
bnt0AJjEfeJ25HUssXTZl948gyZU/rk70/zTzk8vv7CCsePaiWB3H3eeAgOFhPNYRy/geV7dsVyJ
Xp6dhFu4p8AwrKyZTgOCFWpmWDbAjeat47ZFiPWa+WGHSzPRKNNDKVzZRPw6lPKyXBxuJm19PrCn
40YYhlaG9uemsml/QeWdJgWKyxuIPNjpocl3mRhtyEtjq2VlbgpKMNHIw3npLILwrCrIih6XtKDo
vkMLYcDMuNVOCy583gxfz7mQI0ucMhiRA1G/S58Q0o3Y0AXuFlgEfsUVi0FshjShJgzioAUSXpjf
NuV6MK3KUwVYgoZzG6fzM2dyXsH1b4+XK4OIfAxLFURMaXlm6Kq+bAv3FHFGgLHbalfJ74ZvcXC3
f9z/6J33w/cI7bvGj/pUkzxE/VAtfFxsMtSoceR2PF2IgNOGVgWo1KOXg0ZYKefK9kr6WbJkg6GU
ip7N+YXSYjFfjiELG1yEZpJ4dvNRvnb3WoMBNBEIeCyVIH8NaIsHH7d6hAL/yzYUc1nlhm+a5PW+
3Xc/cTKDoQR2IQaW7jkAQWw7t4fi3AsqgUC1gvjqg6z/ncgCh3CGqeQ7L0kY2oIblrTnoxSW9TRb
RLl/t+N1Js1Cc6U/7EkSeYAObFk5BouNTPGQs0omLISHR06kkEhoVq1Fq+hxooPSILTn6WOWAuD6
dWHklQDvA9NHC71oJk+MO3G+vRyh2WVCUmrviJ7oi7lOwCt55YjQ9mPGbckAUeDQ8+rqS03wSh1u
HIq5gJ35Ru/hn7h/U2st0BNyDwtwnhSn4E+nL6ow/im7rWulIE7YqDRvFku9k+qdzQXRIgM4JDL/
jaDOmN57Aan8lJtAvFkFDJbKHzLRjrPyLG1vdBfopMtqhUuQ882yX36vofo/yzzNWilJHnIWXSo3
f09em62op51UYVkNOONZUciGQhQsMjIVhyYVCbqWOxPF/HAv0pJom01PRLuUvb8Ogqo3XwdSfH3I
3DLpRUgrlePqQrfOzjqLhJz67IbFIgM/mwLWNYpk2ztGtEqufF+FkC28LkBx0TV1T6rN54TZismg
dQlvulhj5o0S1JoOEo2YEOzHleTyyOoB6H/XqMyiNjlcSqteRgnmqMz9JZTmQWLgR9kg7fdwl0nh
9O8NZVwvpxuFQae4XYEYnDYssAxCyWH7u4D2EUte+opgZ7a0hs/WTj+OGIz6X8xank1Vc+X6om9P
lqJWWEP8fTb1Uh843LJk06T6M9v1P0UDC7kXWaWjuKgVHEkyV8SOZRdxEfRKDNluOL6mxJ7gDUCX
Mw1sjC6rQxD5BRWCDStr2S6v95/J5zz/G+xihmQjfc625/8snLEsdq4pPFllo+wW2A2mb5BITJar
fTs4NyBpRFG7lEjJC4Fg953v2TU0JGQVe10RUFNHj0ylika2fZZgH4bf/izdogsaOg8aHciV0rK1
EInD0giUe1xKyhSrvPOd7zpLM8qTCzE1TZf6cODwXVbOKpCg7n1fRvQs6dh8EWzx+pF8Jf/CVad2
QlXOZD8qOJ2nmXWd09Zq1LB03Zx3bO51DhRkal+Ae7jNQ96lvfLGaJLmHcQ0LLO+KaJeecBj7bgE
lxCdYEsBv2p4Duf7OpqUOmYl7NaynIZudnPgLOeaxZzExxiSJ/hKzqnskq7ZMkquEYFVRzoYbWUO
D3dteDcMZyBkpK5vx8EJxjAdxOtXAVeyu7RTpiDZhPwW1UbsuA2+KdDuNH8oK/G53I4pA4VMq1+g
bVP7JWAo5nQplZwlZMg8QoPJryWr+oTSYywjoGVgi5AuVRj3GYYEHmWDG9v93dWjUm+6mWmz8fp7
3sEOiyUk65WF5umzWFoTrLgx8CsuJBP2ujVrib6jHEwFBCDShvhlHu34QCMdCxqzNQVtbdimh0M+
Ub1toHbLXDtEXBEOiRj88cBbC4ln2K9Y6t/czlIZJGtWoLVBQwHfj0EhuSjKxxEczZlcpjgPiGam
0b1cF0GG4+/N2ZumWKNlLjPIV/Ea+driaLbi1nfxj0+OEB4flvHEoPH5b8zQDO3vlIg62rR21q4P
ahOdOXIR2hh5bx7Ff6ZeWs/nXuePHgF9FcHvewPupNLj43Qk3DMxCNnqL1LT9kLQNTBXTkW+Xp2u
Z+sdpRr1tvcaVg0DE9eRAQcHIVtmnFBZzjBXMSphJeewKgfUcPXHDEanZ+DWvYqmbSoDug5It2SL
GfBD7Ktq2dCe10YNzkSuHjKjOcsBNuBWAb5fM/n4Rndukn1gWnBEpzloXmijCE3F4/Idl00EdyRq
RuPbaRHe+JCbW7uDWl5oy99ZaARpeF/67sMzY2cU97NZXdZbgLpnbYMA5nF8Cr4VdpIurN9tg28s
fu3QsqiLfoKHea9pT9lJunu5338MWzg2E8wFydBSQirCzjkUXlpmenU1XEbXbRvFxj0u9PWDc8yq
095+cCx3Csb0BrrguWxFEdfprEhPDH+tiSLeUMBz0LX5bHeEDeIGY/1zuHQsuYEtFslbm0iDboQ/
09zfgDhjARIn0w9Snm0d8dR4YU0yg+hbKGdvPKaBuc9SpFVAMrRmwIoj3RXJpwY+fgCAyLqGUQ2t
3QsaKtWXuO/YBtehtHniRsky+R5fPggqvLWPy/ieJ9Q/omywg+UEzssSZQGqe3pdB0/lzwvVW3C5
QRvodUJCiqYJ7/eBw2m/PAYpiRlJRXtUIG+JpNVmMMZ9zp9jw6pChovYzdTdemCz2FEUvoRkzs65
H7A/54pH8uzW1lRbk0Ohz68SPGJEzzYbdwd1VQWtKebsk1tl5jnd561YVLnOKEHAlV6O0VoeH9ES
DZ3+ePZTxEwutgFTKu1cIFN8rQ2hTnYx1hKFV6SF6npNPqLv23DdfrvAvDjUMGddxlRWeOWYsfuM
gMxTXuVZlIeI4/OsZfwQHCfXNi+uZz+bWGf5Dcll9k0wbVejNyky74uTyzxlB/JtyaQfMO7Jv8hi
tnyue/m9grBhH8XYWSjD8pdax540qI6Rc0e2HYzHJkJbi1HmXGhhCzIJF36j6vYO1bxJrt5ZJMzd
4PJOUkbzkjFdsrghYKBPBwQrTuWak+lH1OIYcgCOFuKwreyqmKHSYuyRdXdJAHyYoh35IAQLHXKd
B2bu9j2BEu7qjpNt4h1fp1Zz7xuhjC+15zobJgVyWEUH+EWpF3m/7tGHXBoxhLemelc42HQhAoVm
9vUzTYQ0IONUaVACydYwEWgiiyR3b0ZMNEyaTf147trgxGZ/wP7+On2b1+pLHZq1Qgq+R8XgBcwt
OX8BhISZKYawvQPztjHzjCo154lpwcM5VIprVnkl3X1+VYszEtMbaEPeT1bKhdzu4zjQdO8tGzRt
3tQ24rbZArM501Dy8o/DRZwyIfLy4TPSzUT+lRyG7zIj16Aznq6r6fXCXDkMSsoMySn0k6ZsbuyT
4ySkXSrpb0wzpXavijBqSSfc1GQjQSn05QltXWF3t2mpqMITGANGBzt8whkI9/RQP/bd+FjfnuAj
bvTHK6dSo1APbZy8Fmn0/coAGiChHJcQCTYdk8YqMOKM7ihJSyxwe/Q70PE3fUPYeEi+E3JbJAmP
4T2llkH7FFhDVG8sEZNWgSlOj2IB/t8hZmj9+tgR8tJSp2KhG1f834lklsicsTvLb64iJWg6EiS8
Ju30R9yDmBeQOKfsuo1qpCKJ3Xip2BobVtMKLCH9wOf2FU0DJuddj8inWukbLgKta8fLSuzn8cSb
vdPuHV3tb03yoyupVVMwOzxlOspungiNbrtKuCIEugH8DuaMPcm3lhcXJZ4gIJgpz3l3/12FzVTR
MM00A8eTt/gseXtZb7lUE6D6timXz+NHn8Ho8EORiKBTsU6Pt+iebgaBMTjo5ZRai7dD+z7G77ad
r19xGfcS8D9lSqmVn95xUnsYjc+gVZjqlF93M1iCmFswlFV4ZnRdENZfDkFENdnoV6Ba66uMUct4
wzAVv8cmXTdGVrR4trjb2ioJG7qm//2dtPWdynX6jA6Rah4Oit+/s31pPEA0vQnbOq4FtaUxYWYd
4ilYVXdxDjMqSpszDfNvz2HPzNJJzkqPHCA0OTUlWCoDFTX39ZlofWdkiKWtYVU479bnofBX3qwV
Z8qm23IsmGn/1I0oERx/Hru1t7JVsHxIfL5XfDzVtWUPeLIlFp0skUKQKp+SsO+GeOyAaZz7PNsE
REn32IXtKf8WAnuNeUJSo+f/eSsQWDVLAGL5oLJ2eSMIQHd+5pqH+Oz2uvzfbMj9m0NKLs1dW2/M
CFsP0KxtHyVPrFAbkjeJbva2w/6kKwgaArxksJvJxCUGHxQkrpFitqhzW2QzRw184/hSSjyysMQp
ytI7ANt8YHtx+XYHlHC2C2whCj2aoDhJnvc3H3fOEG29lkygsfwqPIjwH/XJ5nU0eX1scSXC6gZy
56Lhs7X5S2Ri9FTtuembbzMm+QHakOHWzcObRuq99rc2BmaA1D7ue311uIRoIrPFdtUr30IeFd3c
KYLBk2+6ouFJTzbO9a/Ww3BaCXSdHW2xDTJLM0b4WO7+yw9be65m4e5kn9byhBgONtvdZhWD4stP
kFAB8amSfSnK66rEJ0ZirAB1TZp/iOWPOnxZTaX9dPlLHdzgcKhMRRYla3KW8VlDsxGg1YVaM2gu
UDR1+ldASvDvPfxL3XJxmpxymdol3d/qfmeRKKJ/y6Pod+HBGkVF2U47HwHwowBJOf5jb5c/QasA
whCZGK6yRjWuCzwRI5eHnfnPP+JCQBNxMdWYL5zoVtCS2MbQe148GFJMyRC4BonGKoDywPyMGzhr
ZnNm8UtSGv0BuDvvmvkaVoi/wLgd9SsgTwrlGNqW4/nnzG3lbtoWKkf1LEdsxPCgCfSGBt3PRPSO
8FcPigTC2HnT5jbqHp24bH/Vw1FYSe1042mNdSnMbC4/kr9HYbeJ/ZDUjOpOQBm3oNlIrqCR1MSz
DXkUWb+SPAEjPzdD5yjNW8Qq5fJ1sBYqeXjwbQx0kGp/M1/NkDltGjlQFWVvhCyPRsHfU3YyWqHo
FvBElIYqy+j/q1+znDZDRU4czStecLULpJ9M48nAWSCX9EiSJyCtvYhvAmUzIEYyqdpxVjffWNsx
nbGGgP5WuQvFIlPr6fLxudqVT5oX9lyZEVN6TChGoD7+DZ3HDaiNJlin4Y2vl3LOELukaJ501Rew
fz5humWZgEPb5T91ZHzegO3M+Ki6Q0Cxv/7GMnNuHuA5PsMKiAJ4Hmd9EhW484HFmJ+tFguzyR2e
bpio6sWepbXyqEgHlbIXPBRAd6YJk9Pwd2yFde+RhN+pYu32LDBZ6ypEAd2Fzn/T+TKH+4fw5o8E
o8GspM2cYe5dLCxmCfGvB4imbxBK+npF2KFa/aQm4qLCJW7sgeLxZRi8p5PVfU9/Hh31pKE0fSQ3
yeaGJVybOyBxx5rTLeQFLPYxMqiPWUgYRxk+aJIVT6ESr5CqfqYf52a6GZRzpitHgX+fgOAY67FA
eF+nJJ3N98qlaXjrRSN7ay1rZsfAj9rG86bMOS3yNtKn3dtK4FjkGPSOt8Fg27i0dWmlZ0nKSNnV
Fcnh65qxlRV4YyxBYcBcJtaJ4tnHaAyIZkwZQvteX1TwMBJ1Jh6lLZcV0wBioYG68KE5ZeVbknDe
r4F8M0Dtgn7Sr7b11YJz+al/J6uf+u/VVI4opJB5w1CFcZJL2GssHd6uYPJMWWeUXnYvucPNWuQo
lT4J8md6sz7bfwX2Lh+PRRib5HY3zIE7vd9U+cNArRhpNQlLJIyqYUdmjTMJ6Q3j845VR9NKbNRg
soy2ZUMu4loELLn1CdVierZArlJBi5UdYq4eLhbxDBpHnjpxxUBQpoKCUkfX6Sjg4QFxzTXG8CuF
tmkdsljR6rSd8Bu71mZYJGnuFEpP6jZvHx/EFKBa3g2YZXtx5b7pvxiPZm38Ey65WAndvSl104I9
V7nsa8v8ZHDJD2oGkQTh/zJDsEzVkmG6xCMPVPiV7X7HvT7apWtBbZuYt9R5v34KrDuR03Vm0Zzc
TcKB4XjUkdc0bke4f6Y7cjh832a4b3F1/Nu3KaefS0S7DQxeFoYMoyuc6VrMmaEEDDNy4Ewi82rZ
qJTLzgEQZYsesjwE0pmLHqLjUiDkG0MpOLCQenTNMOGktve1YAjX0pCWDznyOXSG/tugz2mIPOF+
MWH525NxdiZJQP32dI2S/lmKu34MuR6doOYPbWm0j8qMVQix/xQXCWd8DcUyeMiIow8evWhQ7AiW
NfXgRfdYof2GozHeYd49gXx8x0LPJFKATMv8V0Rhhb0fwXZB3qejdkGTUazabBPi09H6xTMvkpgi
jWJR8hLZEByZxN/F1YcSJgZGw1guYPpyXEQtMYJgZ0pfbaGx7jdRCcwO7Ry51O8PPpSFKEEsjdOf
jlB1gdD0J/LdugIBgLXDrI88rc1PWg0VkZRoRhM4LZ23cvl2Tqs85ngyfa0Vm9RuYJj0gRiMfxWq
iCDdLehOmEpUIzZG/QibTp0myD2Eamu6izuEC9XqvQcti+mu0T5clYE6tly6u73HUIKMkQH2d4IR
ZjoRXVRMnDSueSEZ4BdpdQtyHnwRPTCKZLG0H4W/DaDELs+seNFvsxkUfJBh+fTfv2yLXxCIlQqZ
ztnjx7FX46eORaUpAdVQdOTUbA+1ULsST2aYr6ukFuFleL33twaIcdHqZad1VTWSiYyAM+bCqURb
U0iuh5LaL/odEdZcdWeFSoBbASe+MMuzOn2326TBH2lVw5wiAzGaQq4rEN4Z/tnplMw4Y0iuXE65
cfGhgu4BAZUYHFqFIH9cmmJEyR4M8bhTnZFyTlxqgB5KppEK37MvQ9yiY2W1AC8b/fkd/TOTIl/u
rWuEjIa4gd7JMDWkDSaIOX34niD+DasXksJOkH9jFunRQwqPNMbE/zGvejgFjEaRiztmWOQpiI/N
fX6AlcqEL4gYfHt1gArAiAm/+Y3Q1yg8/BCqN5G6P03ebSXVThpQgILSaEXcMdoYXOBVLOWlWEpX
DkG1PxwVn/jfu6+lk/OuzbZSUkr9gcoAPt5PJGHBTCGYQetVmEF8KuuPfSUHxJSDjxGckXWgpCc+
6gnD06e6t+l8DLmtE4/kWwh6MkHJSB4yTqO05CGV5up/4CYafaTr22EYpfPQVwZcy8i9a5M3iRfb
kBGq5krey0eUFQwV2B9nCCjXMwt8BNHT6UM4nN/7yNUYgMrwy3+3tO9J9rSZuan1WoShyM/FhnUo
4+xC3S9Do0jfYhwjO/5J8a82knF45fkadTl6Y7vMz+zGyczRtoR2WBsqQ2vgtxfZ1MjfnY9T1UKm
V3lfMlJqnOsW8QKjLicVbQDTik2GA2335tY/da5mm1QkDI/hXxD8siYEswaZEG90UYnzHppw/aVj
4PKaCSbsY3e+6oI0OQrGTihpha2qRGxZbfu5eBP31Stupwfg/4Jdx4+/cWlvOSl8UV7AuQZX1a4t
z3rJuinoaYrU/7BK4SMekmkHtTeaZVNVUun/xZumeM5p6oPqdJRkKr+uoPPCZy4x+jbc4AWghWE8
ZjQd8cyOeIeCJ8q+5rytK2nxSId7FKufAJxf0/KC1AQJj0dh9ZY+EwukZk/hjMopdkLYjUdYt58g
QvlL26tfbGD4OXe1HpuEVKssZZDpEocaFdJa2sUJ/uqWaXs1eMUca8xkGiF0pIKwxMOfYpUYcyNB
wwotDcJCe72EP+R249TH+TPjkFdRkCbupeWalf7Qc3n4awz3oDHb+m802SRGQbFKkbDKHBH3ghiE
2Ree1TOVgayMn64qLLAmIDaaCoDxSYYxEaWUL5g9GlS3YrJV8uXkdrhdVDKtaKH5KyFuS/ZL5J4F
mpqYuF6vqzwvuZZkjwWk1DvjZh6Ua2gX1jaNI/YnxdntF8Im7/bInx8+yAuKJQTZQdr0+es8hxeA
+YpjucJHPZpkGDTeZiPRUJYtHnuoaW6vPVvenLeGJIf+GKtr2Z1KwzIokFBfjU0dGl+hy0NB3gLD
chwEVqh75Og38khMWlzOo0d1hPMZ0ptt50IheiAvaeNraJQFnPbgX3JZYlGdJZT4NbEWhsk5O9qD
cCMoL/fqs5tjrTOSXtNNB5hpmtMwfItkjj0AncfCLjfvVYRDUdhpuK3cwDWYgu5k9n089ubwVf2i
AsuNXmQu3MGpy3k3Z8HkmlZ70EpVEhLjq1ttR3q4UIdBQphxIcdzg8GKcNfP/kILf0sdFsM6BiqY
Su2ZP6yCqf3nBSjHg18nfKWvzKRsxUqRhUPjxYK7K3CLukTxVEhNQp24jxiOqHpIBJqXyUO42MQ5
dMdl5JteLJkLvacKk6URfG21ONKSqeMiJLq5cFw1r3twFW322RBmiISpSOuceIv5vMzKhm4B+Yih
AghpGWSS+uMISQ83ZNDkJ1XGZy/YDxdmgxO9cNET1us7oGTLUag/ptkKHHLK7B3ceKvZii3AJV7R
dSGMGI4g/GypFZHM9l+bZVy8ZS4VzHx227eJTjs9o+rsfgrf2w+SDKYGPRCIfkq6a8wC9q0nrC1N
4oLuUr+Th88mkFsVwT4EQRqbLetHtcRbfGCG/jbKp/xiYy72hGn/R3uP5pLR1grz729pVNWk0BIL
Q3Rcc2eqKQVBkEy/9d7cDYYtKMyMplt35hv92p+itrmZzd6ucREGR/9XeDbk4jc+f7luyu4XE8B1
p5JLGEjYCb9kKP+di1zYd4pgBsTPGnMBNv/t1+/yfCZi7X4MtDb/p7zYMtfgHRW0r9lGUXBBC/6Q
ipuu4JWDQNZ8VLhYWKxDOY/ZRyRTWP9AcZ3hpXHXkDRXa43125gCsWVRTf+FSGG+pWvMhUHKjvPP
46+UPQAL/qwVjyrW2HgQOJwz/9jv0Os6EV/U1Qnw21bvCIsGzV/trmxzilkwOKQzdygWB9Xt4jHO
Xdw+28vlc4QgHXLoxwFioMN0yXeqWdjIcX/SvamkinXo2WnSfDcbs6gPRWXrFFc2qLTULPw8cP8t
F57Qe69WZwyATLzTrYJJPLm/oq2pguOFdSHNaSAOxYQrwRHD3i+KUzz9ftw8U7cSr9KNf3bd/FW+
aGs8tuaF0ZpZuj/hRZUtyqGBQU+DkHJAdDJNjv0RieQ8h9yTIBYMBYT6eB++cOmSdPurLA/R5KB8
8vzGo5cz1lUUdOnwf/l1pCVQf5+fWz+cMA3BrgzSKgQAegRBFVGd43V6Tme+5k4wNrjN0gxkyTUN
0CZIpcPRlSHN8GjYCkTfStWHihjzZ72B1o54P1FRPEmr1BY4r/H76RvxZXEG6L8ppdBnR2UW53lW
OZPcy/Dfme+NYOc0Eazps8ZtH9Whdfqnmmpocm2vuRELtEJuGIcK2Jome+TSDt9dKG6TIYywyvUu
BHpl466pVsGmXekU4YYTee+MxI4KIo3rd21H8Y8dkL0EgyrK5BUvyuM7LzNx5rXqIczj3QTqpr3G
Rd1u3/n1iMAPhSvTrKGkYHKGhenIH9tEqQAxcAt/6LlS7+gCcDA0PaUqPMveXvfbHedpqzjETQCt
saQP1e6aWgQyrQh5aAJ510fZr+KyYLKdSuy9d9KClTt06eWTNAPDGR5A80PVwTZbWzegzhLSN7z5
A0oIsL7pVVvxOQyan/ZDIgQhBphkNi9Cs8DvZBIHoIPj9FMQXBOe+SqgZik0GNxtDSX7ejuSICHI
FNYo9zwz6S/2H/xlL8h4m5RLa0JiQ01a6A+UwoueCsr5lpI0GnJt9Cx8qGK+rHEbkJZ8ba3Mfkc5
7+8dLQZikizHx+kPU40GWqOQamNYTsgpXTVWnC6tvXUpy4LLxKmwlH48uyAC6BpKq0QOeqovlMcK
6i1eHL0ulm8DVZJpN+enBy7HWFd59Hc2IabDQw6LA5MaKpIoQq+mI/M7X68PRvgNTIbCsAET71de
i4aDwFIBTQ8aHvALouTobhkn5n6E0NWGc4sZCH04n5rfWWETONnT9ccbcWMysszn/vj5cIoJ5AFc
HaYYuulpbXUE/bCaji19wLoXq7RLqAEN8sVWziB/imcoc9jSVklMhF33T6YBOJ6Nkx02D8tEYhXd
OwVERaoEOEyAb8Eqh9D0Hb34iFqjB6K1Vh54h5CzEmG4qIh7XiDrVbvs3ZVT3jEwljRPP4zpib/2
qK/OYRqVzRf+5mDIjE0CrLrDEHe96a3BHKdZZJ+rspQ3WxTf0IDWHdCiy2P3WaVemRW6/vUR/AZL
CM5pym0gYLxugGwp+aXfzrn5Z28uGaeTdACkhXfsag27JoBR4ERBCJbsrU+oMKMYCtIbu5fMde2u
6htqEyZEKz3M4wa45AU3oyUmhmKk8zAECOIJ7C9L4GWSrWOcOx6TsAFm6Q3rVSc/RT0qXAhXdRf2
tY9MT7jG1FFdjssKN+suB+pc+mUWO9IzhA9ftOKo0bm0uoIVZOPgwZlCEdQA8ouvrBhbNRhlNdji
NMzTKXePlqRr6I+bnPqdxde12lJ/RV2Vn3H2f1a2jl5OcIVAnI/s0UiAVXB76xe45rvoJMOw0A1D
STvI0rgR77efuihsSnl4XgbP7A2D5KU4hRVRLTmdzkF9an4sN1fNkcXdUJzeCVrB+VaPdbDx1PQD
4zURfL/hrqaj42T2yPogYCEDVb4x38yRun38ivxIorrHegCt2gRRIV+z5vXOHC2kc25i1jDOcE1h
qSqfCb6fBMdKF8og5q5BZD2j0MOjYjIpnP65JwcdraDGjCk4ulO0yparDtD0Y+rB7zq0Vs3VEj1n
vE9VePVpw13OUo5fvk9vmZIzVM4FLe1YBO8tY+MlWXJ4rKGeTZ/rrUv100t2eAmQDZquV6wMqIxD
LvFcA2hrQfLDabNklPaxK2r0HE7nmulQRMCe6ohSfTeH4SNKzPPS+VZjFHBrRtD7eb1E4nqm0iT3
QDQmgTms2y3k5xvJg/bU/Tag9ZKJDIz0E0yqa1VyYh5mnu/RUbRRaUnIuelDNAfbM2GfgBDNpVQS
+8+ivUtBgOD0smMITIG4sLK7oly1pMTPpcIDIwHSee+uNBiDIm9PK2nwiuXgRAOZ6VvrVZ+PBy8j
90bdhO6jDZz25FlHUD8/UKfj9+MqoY6yaiBEr4AY4o46psIs1PaFUw0SXIRxGq5/Z8gMc0SAr+95
LBWs+sfMl1Yj4w3KcUqkdFbU+5umsdIwpXZAdZ9GAYVyEwZy7QaptzYd1Jy+YyAggrgB6WdvLhMa
Iouc7mVpDT1JPm7ReW3C0GffZVVHJ7lPUbJhhQdFvRmcNA/1sipRiQ66Bd2URW6En6K5yoJ+H0GZ
547KBO3oFwVD7XFPA+du9cj083VboTIQ9bVU+JFOeVMU4kZvTU+8ZG1iEruet0/NI607AOSLUJv4
6wqduRArz9tvyns9R6u5H03k73gCH+jdgX5a1kVAl/DHq3rlUmQAz4DSLEe/D3CUy6x3wSJIVuV2
Ek3/OVgA9S4DVqhWdlqB4ebrKIztxuiPg8znP7YZkSsf7ZKHyw7Kc+/ypM8D1mWYKuF03Uc4F3Mo
im74r6MAj7EjOFvvxr16wMrb3KF8tnvviIFl6M9NVStFTkW3+vlM6GICMyNlOcsPLipIDuZn+sUx
mAY5VFN9HhtZmBVpHXhQvpGz6YZa22F9YTzuckQ0V5sIedjyA+huTYGGP3oZ1pwmd+HOciXcPQiN
RcjJRgPZeGfFc4X7vdiivyt22JFn7xMbMKlR45knvogArY7UET+Gw+pTFyoZFZrx6oKtaVWryLJG
UeHKOgQgymXlKDuDQXUvJLo7yijJZkHZO2Sk1CB+l3TkflI/0JFsFCrdi9d/UozNINLiXh+erWWj
HPUjcZBXEkFUQQrHJLlXG++wMmKKFJErWMFrmXEgfWMdWVl3Qug/l0D77oNO08V258Ux82crCZYG
o6wDaNzK8JmN1FH+U+CXcCWOZ/rgo1Ai4H52c2UtuRHkaB9Xylg32KDWasVuOoAD3I6NPYT+nZ6Z
DnQsZq90RdsTEJsFi3QQTZJJRp32TSqh+UC3Aat7k8DlOjc1olajtklPNrLiFEwGFPFIwpfftlhQ
W2wswYfUjlW5yIY06caA7KrK+je6ysP48EaecW0PjdxXK2mQelpYQIBZhcvldnc+dDFXlcq0tgRP
qoH54giyIKQW9jpGfID6ogJvA3CbPW3YeM6GBBYeUih80bbTCYFpcH80MaXrWz7i/b7cIqfttqwH
d90BWx6gERSRiJlScE6m4Fao9du05FzzlgOvphC1UMJ3deKKcFKOBzlNT288LNo7bwDhKrNJIC08
/Sm8ykDjPWn1us8LZiEShD5D29D2ID1tb4HGGLdaFl3cvBhU3bbNkiHdD15rZHdV4STqvX44D2xc
WxadSSMPWMZozN+hKXjoXxn1RtrynqamwKiSZYF1uxZSomw7OpzwkBxPSxy1J3FGASgPlM/x6B6R
MRa3kA4VaCq6O69lsp+jdXsjAfHcRsKMmpVkR0jGVIw924Pg90l2OK0wNFdYADSJL91pBF9R96zP
6fPJL+8mGbh/EgKlcNlpKxZCnWKwh+E+ZX66KxYDXnzwZx/B3AU8JDYz8zjtg+KgagxvP4JaTn5s
pG39UnaxQwJXvr01D5oWBaDodvXtBxef1T6EnRSTg95/UGfsdO/EPY+NxNnVNNH7k4fAOea0d/ua
iOTkURawnhphJMxLPLescka/FF3Onv9lNkgbBq8xas6fvFnyY1TeZGxPo5Jb+Ta873Ckig6RDy3H
kqKXykcUALjnD5wLNOIluaA4bEBJGyTTb5ONi4KMxylJwVmEc0Zjmm1mswF3P+niCxFkAc31PB9A
Ps+Brq2XFQ+IFRlQHhNeRx5Ym+saqYxAhUNye2TyadLKJumEQbjFTZo6kWn+As9Xqi1YVcecw6/E
PmUjHyVxSZP0wm06RsotplguLeoPYQmllehcjqBiSXiwcA7dAySDJ6oPl9a0m0XD9x9nDraAOXu6
0xGUFsiyOht4083ZiJfSXXAmXCgFlwiBgW1g3OaJJ9TmfQC6nbFnZwY+7+9PM5/7fWUO+YUDSQ7/
TZUHVN8r3/pUPkgx6UeNkK7E8IMDfsn11PZvkXvk3EW5HuYlhW4fvAbFOz7wFQcd/CDId7bQ0X01
l2de10/hdd38fnUV2Izf7Nrvp3SAJIvvR7FxIopqRnarhZlurQLf0LZSFWo4+lm0J/QcmUtagYPH
oLJthCR2qwGZGWrGg9g5xKfpsX2mF2AuLybY3x/REm/agFXdEEQPit3AALN3x8NlbnGm1CAOnd70
kO25T+erVFTqMCgayB9LAVvSKxOeeC3qkz7F2z02ujjYMg8fzgsLuOVYCFHr3Gt1VERMkfp0zjKo
xOOggezebQAlUxqjPwR142GRVezpfdqdmovdNsC4Umh5UJpeQWL8HG4079B3yA3HxiOoSsWoOMnS
4Gedmn0D/hnotIlX8XRV0+MPdeXDi3CYKx/wdhiQ19VwAJLCZsmt+P2A8AhgZmiAljZWTREy1OXp
OpNnHVllzIU0XC0Qd+Tck+W4yKa2atidtcR3HylSHwJGkv3bGl5KCWvH72ykt0oZrlJLgJE5Mo5+
5bMeu9sUYTv0gDGKYo/0lRTi3vXrVluddtuwzIb8NLS3eF6VhxgRi7qaAM3tfJFIMng//+3CrGo7
y752dzZlweJA4e6H2l4vFgz64CcLYsnk3zuxGwwftt3Euz0cVXCG3HJ+wKOiyZnV9AYdi84MIOA7
CISfVbjJqgytysJwjoza/mfmcIx3bTMqAhXKIQ62KdMOi7jXPMO2QiPosCtTx8xZ7FbovKsKXIlg
vd4zNtAbXZGVL6f9kmRA1YgXKYmVmJ/vdS+jM35y0tqV6AIgVSCl3tC3YQIod+ewnm2KLW/v6vds
7zCxmEI78E0fNDk/uSjI1tIQndPOsoItvzLSpQm/hMi90P0ynFkmgFJ7Fo2On37pYTyb8lEJqGtt
CCzBMT1MqEr04t22uHXErfleQpMfK7iUXO8b00I8bpPm3hU/hd22XaHQ/M6sfH7hFJnZYaLzbtP/
OmOr6YW6SST9cTSqeP4drqu5Gbf7/6GaoRclhyastEvlVcYqOAPZ/uc0xsh6mF5UYHF0S0HLX5yr
qyzHsy5Cso8hIf0Q8yBlvemV4xauAmwA8Fpec6mSqbx+w+NgmjurCe2kYGPhVeP0UeBOb8gRmFPB
77j2LPzC8Df52fK9q6m9vC8z/oer5BEOYq7bqjKl9QiE6kg0eO3KUuUN7YBLO6xz/McJUyF1rM5h
tPQeXNUJlUWSN1A+IH5wiHrnkwUX9I1QMVyuBFaiLV3OSDHsJyF1vijAv+M8z8VNCJWd6IVuwsla
JFJquYZMn/7Og3rdeFgXNeO4Om8zxtdUoTdKy+xFTaVgeV62HawukIEkMWq/+OUuiOWbaVVQlCOe
RkEqUEub/Qf2tGXIWh57sF01lTJXp0Wnl5cSAX0ZtFB+auWKhzIdnHOiyiTfwAKzhFFeuMSjleyV
dL8wYnf87oxhVHlit4NMvlpkDUpwv+fb76HPNYBXIx30wB1ehuj1JmotYGPaSQgHbMgSpXY3neGj
0e3I1+S66KUUFQSRXMPIsR+lh/61PwVAQlyDFcx6oUMINEU0kDK8giiWy5AH5ow6M4U2e+l9cKRj
Kvkxo2038EDRBQi83JeMEEC0bI6Wmk4DGOpHtSs7R23jasqhfHfVpfnuhgalC/e20ION3+SnzMLz
3jRL2EE6YSuUdwOxkAjojtmL1fDADkBBD+DF4bxHJToBVsbHKWZAbKdEzPjbylHLaOK6zMOngzXo
+OsPvFg/gkjKOXgeo3JB7hylQUXNwt1OcZJf+7cH3IlAhn2Skl9FrPKugshjue4YGE9koLq2hFdK
h0C95/ziWsFPKThKtADQ2rlUM20Bkp9+MdpmlSFD0sw6DBDsVjQ3hPZ1i4NR6e7XEBbkZaeot+pI
0LHDS/oqd5o/g1zzWQCJ5RzCwJ4FyqXgxwPNDQzpsGe2x4Xifjeu2VGD4FdhIErzohZ1rdC6Q9Tf
s7mOJ+/RvtVJkN+lLh33K9f+4483QIju7WLZlYqtJ4RiRkwaJFlgGKIMqz3lF/YC1ICNpnSInqMF
PN/eVX1xQBOnmCrK0u0ArFHkFCqjF/2OUY7zCvU5+aYfSCyzK9Z4cn5qZ+CvQ1JLYMSvxDzzs9IB
whpNoudwXq+u43s9XNHnatqkqtj/UsNT1E18WPcX82q9fHdg5bOrvg3gGbkN1gKE8WczrdhApsf6
nFmKtAyTeHOjo3oiK3RpR6Dk0uovhfd8hfi0Lw4PTB8Wmg2CFLi7Fbgj3h9lByjZh+epljJhV0zM
RTC3vg7NHB5j+HeeaoeGQdWdezBZVBs+7jE/MSbJyN/H9dw7te3tJ2vqpbB6kA2MU6eFCzZhRDQo
G0d0Ti/xs2310hkUvgtINVLP2ERgukWRTlfiKBgSZ9OnT2gxHTxIagSLz/4rnDOZHAQeFixhUABN
F/aSgKHo0bq/LEYjItqR1vkSq26kr90LioCAVv+LNlusMLBGWNaarw3uy0xz6w4eOgbBvIoUCXHv
GEyG7ADSPNzBNHoTi6nhIxVhQihPNH0d8rWws0G/e1ReuIQhFo9dQOIB7MklBNflxpgbdXRTT3p6
R+oGTqUQvLDgsc1U7jvFlykS+svY1S3aC1CrQZRe11leefkLiBSO1FokbpyRkDNE+LfiPEChVwL0
EKai715TBMBgN1J4zpy9KPFCz4xoRlc+XtoyAittBAZJcmTPFx1ukgtFTmWluWahr7HKfyeAX/ka
UaONldnOSFOnCS8GTmYHtUNuXB3LInw0i8k2/HlaLOOHcuIyU0GATo+ZFesQwqSO/Yitc8eXTKIq
GXxi8R80KNRWjI7zJA/l1KkPUV07B25B5ChKaGJGUlvQZ1fFvB6Wpw9ieWCTrHC9/QOx7SK6IfuO
8WNJv9lTuLQe0Sun/KUCvreANqYCMPCfvL2mjqlKab5OVhxnvUmsgOBYTTeip0PwmEXeHsmNoPLR
BRfWSCNgME4+/k+9nM4pI4ByV8DFFEPB3aR/QhHRG7nQo+Me5RXR4/NVjQMRsqq1jw76DTYnaJvN
iUfyKMXPnCtS4z1gObeum7ZEqbxZo83btnyXYWaAZvnJryAEk6UpIBWvWtW7DJfD93bxWbwdNWTc
0EJdwE1+O0SPXIgXjdmEl9pCUa7KViCEJxSxp9EowtUsnBrq88kLgp2t2bmsJwt4SjHs3zugN0Vz
OyGW+xs/q+xm9GGEJ3F7NK+8mwbYDHo7EKxxn2f5wpSsUMOGqqo6b+5LJb+5gwvaluemIWg7zLzq
kh6G/Pcgmdr4quwuPfwURtHUwk+mkr97SCVy9oMemNB06WukGEQutcyZSLLYlKQXGmPYbqvIKvmd
LJx5RwD1i5iJCuxBD3OXmT9qq7p/thOFhGhqQHlFDX8ZusNwe4JZA4qcOxaKHT7QKSfqX6bFB07p
meEnF8wlTa7/lK3xkWBPMFLWQiOui4uzwYpeVESuzQdgDfk8vts3PSQXlIMvZw8pfqHTn1vWOT5W
KhgTpzSD+LKoHca9DmZ2Yz1+jXZ3pb7wruOolrchZMyXIbdk/7mVon2RuBZWDBYP+VECT3enGo3B
sfFmfJKp+fWIhe2XDLVBf1V7ILo4eVc0byFnuasxQcACBFzRjEh7PcJ2U7USN+IpYQhWdNYCqmuz
4In4xguG/IJKn3G2r35RuEDdjlbircB6hxXmQTRzf/RBSYBaobqZ8NTONPUbOe94NUtDsO/+LHqn
gARlD+YbvSP1geqHck+ERszy1dieZXEsay9pE7db908K8Uwnk+0JTUzXK3FLpqC2CEwzZpRQTd6H
JjRmLIBE2Pb6l+PPEYpcX4xjExkJAClHEzDEziLrhlO+60lcnI+/KYEtk8Q+FPTPjR7Cxe/JILj0
wdEH39oFoxATNAYJh7MBir2uIUESxtYF0dQ7Tjq0aCBXYxDIa6h3A0bUDEeEm5QQl+PYkouftAhf
3UJfE2DJ9OPCtZrBlU/AxBD106QVlRrBxogyO9N2Syy5scoV3GGZX5l6Vv60MTy4TgIYEbmBUoGP
PGwuHy80RBhGfUceH1D/hsazTWnMN4Og8EtYcm1Z93H3oJzRwqIoAn3sZvRUdCOviMUNU7HSkl60
tEQfJYZpaBgZ/IV+weDUJxfH7Qk+Jc5hV6U8ob1xBC2Qmghg/ZPwe67RktO5JI3T9Td5IIucyAAM
Woe67ax2t88zK5Xz0mivv6ze4QxEWzYLZiy7thlcsyW6BzEKugJZmP5svcVcVRJirHpTfbiF/zis
i1yMfNqjwQJ1R8NOGIHo4uceLcleoXfKCUDe1SUVVJz1267QsucORR4TSy2byvU6I5XAWLrEYrgH
8nVFEUyMJtDn1DE1U5+mCGa6eE8m76UvRNC6U7Jfjhn2U2eKTA0tVBKIYp9561H8dhvJF0HPz0PI
z5aE8apqTPQz13GZg3bTAuWqPnr9Sf3iJCrXaddpwvuDxQoUH2DAZw7v9C+LSbxd7sXsMRw3moIz
PYnBqypRAmFUJ7LrAKXc7iWkYrW0l8ZG8249/UiULfx4lOLs1OxnXl8I2lLH2beLilcw2f9IcRFc
x4Wx+0rn5z6zdI8ajYvMGiZ9A+fZk1qp4i2blq9VXzu9yKQWXVEubE5K2DPdTObSAG/x/ww6rxLX
s5Ts/Xc+VbVjbJW1f3pItIS1Uym7IBxx+o+18Ta87kHYH+a9ozQueTsAthe4gXZsh+NDC5SblGRE
AxrvFACGeJBU05ZyHZTbMzQNuQqVV8ZMxELpDHQ41UCXIG61rirP/hkd4MSFps9a2SIl6h0XafWN
swJHBoCRHOFn4F5vfSzLoYvp9jMC75/xIRgmahD4CPzGrfny+/ntTQ+zS2tek9OwF4Biz91+peoD
kwnR9xbYChNGloO7c4vQxKxwuV4BIKqvWD3Tiu4w2fO3wu6BVZOJsf1gjLDCiB65+Hjx2NLo2Q9z
NQpROBxMLzlXuu+S7DWnfUe8s8mnMzjYjdAXyGcFhG1ym4bGPyWxIXVsyFTIdURSr76IpcPcW9Ag
iqA5J1QLTodnGnNgGwQI0Z2hFXdXd+y026FnyGyrjnxzF5W1pF8veOH+Be8fUIwP/KOacqurbNwz
rCXIx5c3f8oiZZZuDFo+BkC6lNEdXkluFl3ft6lyBiLY/r/hOOd03C08xGKLcn/lfkOuGxdGd2Un
k1c1JYxkEVGf1WworsnIJvGYmklT64XprP7KGkOjX37gh98UtMTFGgCkyXxl0gmzA30jiTcWy2Kv
bZDYXNeAUUAEeUZkX56kgQ82Q8mrhAVKJwqoRErInTkwMvP6sHhYUc9ljdM+UowqIviZR/zmMnHv
96Y6um8L+6BVf3617HGx51OWFpYZ3rJGTa63etuKXPPRGpVFeK29NAYMqcnUpqEnSrQ+d/bZGbum
GjfLVaiEiMNjwWzFOCZj7No9nR77y4eaN/IDE06jnu2NP5X/ZMbad6W48Xez3KZU5wE9zjCECW90
Vg03UGHZjIb8AuBKtgpwtjdjtpRwTZwvnt/Mf9hrKs2GU1nvPS5jV/sNBBgASY/RdmOluDats+bY
/58UPcCqr7Tq6M0zzGDy6LtR9XGIO+vT3ACcQ3yOhnEPaaCfCZhCUJ0EMy4Q6JJuv7JW4Lqu8ri2
Jst6NeoUqdyHgzY+cqiQTbWYZ2TWdqnCaEQGJB/eKHKgeLSGHwwiaHYGCrQGUJIv0sOtU9TWM/Rd
iIBAy4ZLkA+4KKwPs95PGAQEW1NcQokF/oJB0o821J7yu8hh3F6frKDZPuX6U1slSgYtuAZ6+kZW
P2qX6lonVd7f+lu1t38W8YY50Q4hm9NH8L1GSaXOtcT5uan9e6vAOKjMrG4vKXEpREQryC7xon/9
YuJjGOFjg1ZYhoQxbf7df2O1yAJXKY0gB7yqC2H5n+CjiQ/NlQF95rtdIijru+LTf6ybdfa8Y5ki
A9qcV+t6jqIKYkXu+IzIEb8qtJKipdoRHG4Fy0SYwUMVV4DEp4Ujc0FHg95Sf6+aLmKwX05a8XiB
lTaM/kuD7fRfQjeJCclY7VEy4zIkJ0nPmkgBp/UtdGNARhugdFLlwAYQoYrkvoUeEmgaVXm2wrjO
VC2aup3IBXUWmdRO2DkdA8uqLGlKX6jY25RmXZPZnRs+alecoPJZjSsEXuA7eiqyvU3CRAPLOPwf
NGg7UswfLmzSuVrEJvRmSVLaT0UFxfjJdFvv/2FYGDYJCz0lb6jgB+s3dyHOokTPhYZ3sxnzvWTe
oNZS17gHm99CpccFCEdjjsZjRgOAJDhYmFkBLOFjuwRAhmaXiAXQBzQhQVOD3/bnlm6raKOx+29B
i2XX3JUqDMwOl2t2FHt/24FBrM0aA+KXTCFpxhjNwPHGZ/DA5Requk/KHUb/2p62LQGkSaIYBCCT
NIqGrJkCGETHQZRc3ediaa8j1H7qjqBI3pLnOiMUYkLVYaourgu3TOiEPNUkpVEIieebgKBHtDa/
R6BxeM75U6dPnKRoZpVA76UDjvz4U+fwudjxYiL/x7LZr12+rPx5omQxi6Q6Vyr4fbElV2zis0Fl
k+1VWFXt0RW+p4U7sMNQrbkCLWPTijAdwV1NNHcbeaqUg/lTbFgWtFwsu+oIGDYfpm+3ogWTar2q
ph4zN2syPGIC0p784b97TeIJg46Wk3sgRzgVGMUxsoSMxDctLcPoUp27ZJg+lfvJCry9QUS2F1aL
Fuuh2tVEuoRMcfWyYhpcPd1TLQYoekysto9RkGUTJ8xUOtMiySy+908w1rvt8JSkRokVoHM3TxCy
gCZhLLnRT1D7l1M9X4ct1K/3hBFhW1JLRwmrPivy7Xp//FS3P3hRpszQjPoKKghLa1OrRI5VevS5
vLzz41LUaMNsSU+ZjIx719L5SSyewp3yn0xAotwy3LET+Wf7Or1gazeGY8sQKSWNSpNDr/gQp+u1
DW1/HMVwjTmCA+yZPtCyMEhoQL3pr7sEZyfIt+kXqIciMOQIPbcHuQ3mKZan6TnjcRchDenW39x5
2cdu1AfTN16GvbQKv2aeEh1JodQZJDlgJlZZzVNpC4t6fCaLjkzarSqsG2vmjQA2whzf1gPT6QsF
C/d5WoPBViPru5ZSDhLx0jD80PSNMSRRzo8U6t1kC0IfE+TwbdMgD7fY1PfYHVOBcxNtlo7LJR6l
d5MwZrrqkk19bkw1t99TLL4eoOOAppgLgIg34gvZZAp/eBLkpcfwppBlbVGYoVWJ1CrVL8GoZqTt
m56ee1M3js9UaMNxWTuFeWtIwvf9/EXGB5g9Uz3b8h5WWfFmNSeHHjLoIBGO90T2Mw7LYP1UCBqD
dEVU3HabMCDcg73z40l+8dTo1lp5CjxbGrkdgHEA4ndNMspbIrFr3QjHrrctIN/AjhUgRmS6xYLe
ueu2TBA5lkcLI6bpwQFceX2ak+MsERnX2vbMSmLF2HqbphZUB+bjBkzbdoAiEqaNEtXk+5FIHkPg
sAnKi2pbcl15qPUvPX993kjOke6jO38vPd0b45w8Ks6fzxXq37/Msy45LC4vPm97+6T72cFFkauX
vZLtPaMDvFtdko5gUYzIfcPOQeb/RPOqbvzjtm5DWQnnkeMhod7jvXEbESqnhucOF5YHSomhNMlS
FH90VD2EU3pDsf09BRGZQztnrlxsb+1WOxwsx+g/kx92q95h66MMigmqHTruTirqWjtHHJSt8vmh
NCUdQWpadn7xqlevm6dGEUp3dfnNYSpAopje5USMlebSLcGOrowuhqEQNWd5gFV255J+M16S8jny
1kMtYpeHjc6gEKDwJqtAU1HkfyhfyYGS13ntALw4/ZYRtnWP178AOMybr0gxVh8o8HqlZ9BshMDo
STsWO97KnzLhiI0dZMAa1nnBUbtjnOVT7/KlPX3RxDIH77hLbLnCz2ireT59Kz/SjPJ13Y5X60ab
lsHcQ984BjFgqFejU8YH56xmkUn5dRHFO4cmHEdd53m62gEMsQoPxfAeXtR1WyHaEz1FCfYwZ4MY
u8YAzgvPp8Boc2qJmuFFiJ/FAMkg/OBHn5hsnj+qSDW7YOpyJqSmzRt8A7UvN6E5HUoJCpqi6aBL
aNfo4eLvPSd7eY2pNKRFJhL5SrohLyIRtgJ0zNyctrnADT/fOGdwyf23/+4nE3i+7PQLAvP1rpje
iZF0JNdgyAEWXroHGn1gVKR3ys6xmhI2kxKodRCLxdqWPj0QHP6ywOLKXXYIRgA550Ib2uA1edEw
ufzS2en7jeQWiJGwEIlT33e/qw20vObSFautTjPMpp5HNhXUDCB36zji5A5xiXTcd0lek+PCHxw9
ZUseqWmsK9ranDjdEV/1I0Vr2AfdNqkXm+sPe+Xj6Ro1XEtfPTalJnssol0NSZOF3KPkQM1gv8AP
gui6Q33rQ2f/N4dc1V4xUY5mz0DXSsF0xORb/t91lZoe+so+SZj4DX/+44aRxYa1KLyR01VAV25f
2NA7w2GXXxzd/n536B6n/o+x9tbAZO75XWUsHQgaTpQcEQMZGVurhPgywKa8qbEjyJ7u5bzxk1HS
Q/lCecPlH98BzAhiIB3XzTMffmcxG83rx/Wd1LmlWFaBrCi4NI+A9dSe6JRmVv9ILBCTo8WeTp/e
69euL8+WpjbMSztGX+4te6Vhrhg2meOeQPrsiPCRYZvf4DOnbeuX9Bo9nnnl33yaO4buVrz8TkMa
oRKx4Je6HHps9KlSQr88sJmoWUjJ6gxIoprlxY4ISt9SWuzK4CDI1aocLscOhcCwQNsZAe+bieoT
y9wBpE/CepyBBTkuRVLg2KYeNDdqLqThEGvcFcZ/IA3LgzUgKKMthN7ZDhv7yaMh8QfhJXnT7kCQ
TXVm9ehFwHxg5YgUwxvP5VKb3K+9vYQQfrR9PrqBX7VbXTdHwMMI+rqbWITJoPlZZDk53TJcGZ+D
9UoY1u8wPOOQm/ugFO0kE/dHxKRQmmwyVAGYlK6gwQ7JylMlrufTmo0jZByWalw1CWifXUCrF7zU
8TI7LGtiUxL7zTsCu47CErXu/uZ1lQL34Io2gcmQ2uXHL5+ipDEKtZHBFDpp6nTXr1GZB69oSPhE
NU4I22KSLIymCYGgcGo8PLaXO5Bj7zu2+OoL+x1KY075UDzyLJb/Ai6FpIt21RzRw+cHt4MMSD7b
kM52Dm2iBuS1DopYx6COPKGQmgNoLj91hXFqzQAi1B1XJ2sPVKutrtTJNq8Yi9tIGREKcS5sgU9y
WgjIa7bAp+AL+iHHIPB+xm67aqok70PdY/QiRvLfoLTk2mycipTNAmakGkzjn/FTYLSZPKYY2Ud0
Ro8YoZT9ylv34TN/hgVmiUzFP5FSNAwQnIRPV+Gqjtf3uTa/uhMiovqwj4AjKB8l4u7eUz91uHiL
81ui7sH7y95RySWQu2K9b4WWe3kkurryhChjisqAePI4MD0zTSmk+QmHDo5uQYeQt1kh8JjlAMnx
zWjYS2Ihu9hf44NjMIEnnjR2idpJyAKCJuBfJHk0vStMZ12i6bs58/E8VcWpdd6Fs8GkV5qxf+o6
R6XuB6tsTIlnLa1wgMWvmwdPL5XISIPATUWGljPs9SruaG+JOl0W31PMD5zJTviz5Y4gYtArc+mM
ghDQ2GoI68s5Ljph79UGnUaN1VtC9wG4HsCJ8NObaZLKQQo5ZxETH+nN7upVTNgMVY1pB0IHAt/l
t5NlU5X7YT/syP6EoeST03IIU0Mc8pUFr28wYFHLkkht7FTwTBf8KMKZj+JylCABpF4Wr7m8islc
4xQJyiKInPb8gB3MwRboGA40p+zWJWsiRITzGbh87TjCESZzvJEjHNAw66vtOQfrgzJxQWcUpwIc
DopRyEfKuyE8Ix20N7XQM+MjYbnY/BAStoDmAZHgRb1qfBKz2Zr+tp8pcfndAU6L/XOz5Xg1VKFL
kd4X93V+CztL2bO2JW2CjvOnJZo7cAycbMArUdxZNg62wuadDTBgOkwhdqig/6xfkSrU22h+Yicm
727Q8rNHvLVFCkbkt0AlPNbC2djJ6nkLw8Go6v11+kJJT4g59OesHDICucwcNKAayk9PXLOdC7SW
G2nVA2yrGrLwbn2NW8e6SIslP11cK0sL3OBixhq+jPF7mdaoWKDcWw+5W2+3gxJVlCiWAk5l3qAV
U0kmMKbxMYxDr+tvJgZ2L5iTIMuieNFbtt2UUHfGBN/1kAOUwXbIyhUvvamgjOxN0hC+9erUoBNH
/ZbVRrjJOJcChUpW9QPsOvM8wbeG/bCe/j/2G2YbJiRkq9eLmYP3NVAiFF5baXH8vUNM4v70frr5
S2xjm80ybyPNHq8dPBg8DJF4zJHA6MRUU0p0uViTsbwue49PQJ++jcWM3JSQA5rc5JlekYlsKXtz
QDHJvsK3PA0L4n+z51O00ss7jooovZE3DEReU9JiKLajPOB1xkVELlDfyce45rQFEBurfYdb6agO
Zu2cbs+s0zwXqjY7A3eggy25ANMKyNCG7TO/AgTq+kSb/TXqUOwga/mwYiRy4OXM250mELW73smT
h214wTWU8Pccqsj8zxsDCCmIGI8cv7UCYySEi351zYuuOjlYOAQEOuR9wgO1c2PQ4nBrEa+Dlp/3
bJKWMvAiI1T2Ned832ZVoN1t/rDlvvjgbJJUaOTd08Wpu3m7eQq6kvsvLwAdQm2BSGhbVkPgEwln
f4FDdfo3uLZRtTFfMHYzpkOmn3hHTI+dQi+SYmhgthNU1bXocnG2DXxtTTmOfZXAhocDxQQdjeNZ
uG7WbA6p+fLFP969EoY9yqnAhQKX7S3WtCumAqpilYpbSX2uMpnl5SZV2hWeOKc4/vBU0N/azB5l
L510dgnT7knAhSnjn6hQTKR1w3CR/CGSlqAsw2i95xJhYyd0QqRpcRDOD8pb4Mh04TOxqlTChr6O
uCPV7hDPqTQ2A42yUHpA7bFh6cL/tJbSkRssrrQ6B5GJZy3y6ncUJ9gabxRchRu8na9/Ny8zI3SA
xaYQTkRRZaZKVo/x4VNT3PtbwrQa+xEbFeg3JuWtC1oK7RNQV9sIuX0+3iW0B7T8vZS5W/e+cmQ9
P2Oe3Qoh4NF67PEITn9VC0a4Xra8uVzC4M6EfLjUt+daZdkCcYYHR+vXWymYT/x7aDvP505Fdlt0
4ml1mKVeVe2LFHgCKsEhbmqBXi9NtirGJnTJol3up9RKgmgtGMMcUhgKLhJy1rqL3QlfP9/K4zvD
nR5hKGFwHEOE2IbTM4HWrlm0nK+TQn+zkO52E/lb5902Zd7jdIleU9AY6zCDU0RaYrSpNkRzCCru
t+KA7+fvI2/BWxYb6XPfJ4TJ6ElIqznl6Pr4oy0A97T+zeuUNc1FrnUdiHAU8A3DrK4ElBzKYVZg
MeNb0SzP3Ascq2NyILDJ/adaRZeZ2vUPiANQ9pLnBirQg/fqHYhQkwhtngClsRNEyGh7iBifuHvu
UOR2lYfIq1gPIseV0iaVMOi5Ht/VFrL97QU57rFU/7cJn8+90ZzEvWQ6AmHWdwc3aCteCFNa6JLa
iTWyUZd1akeS1bwheiW1d2eJAb0jZnUOYH04Dhift9pD01ZBJYOu/NnvQZTpOOQhjlc1zSZzqKy8
Neodkj8mxGQQzOas3YYu88ZRwVUWQY14vGkWgBnCf4cxpB92NQPSvp+JgwCylMJ5cfDf9oavyOiY
jHet6eDKirFMXCMtHFP5Z63v71AoLXlnxE3MbYirejxjKJjF1yOFaiVHIMlZjD7/sQ7JItbm3uMG
bHVNrQzhB2UyqADDMcipMHvrZNMv6lSmdWSXt2Vwi/uSsYVwc49HAoqz85mPvXmISOacoxwJl+x7
JQk0CxAcv/QlU4WOsuSwoGmwBbywVgNm8RU9pJd4ebz5FCkdIqnOZms30PEmonIR4fEf3reHBcM4
0RqZP+hti5FUP4HT0kfyQpYE5jwBHKxLyKWZuxIDxB0JcW/nL5qtJrHFTOoZYyIpLHLmkvq5vUMt
tmRyQGykZyDKb6wCexqSi2/z1dK2B56xym0HhtuOZta7jngQDU0gz6yfre5VtpESwNaBlc8BbQhj
5MmUHiRMiM6pl7qQxS5zeprvgQ8zvERc/cwTj88ROkj+u/3FwnunrnUk0zYxU7tAm4x7Bggr3mG8
kGL7GzBAzuZ1X8zTzrMjlnXhiKYCQamDVuYyrsE2wa3sb1l3IFiboMJ60zLnytZGndgsvucbKap7
cjdnJN3uMI44hPO5FGdEtVPdVzUOE36bvuQRp0i+ER/6A5oxxEA5vpz/IP5EkROHIhAqTmjg8K6M
r0B0sR8a9FwvIc7ixsYFRM/38j73DIv2jToOtOWmq9s2KeSR0BQgIdj78T7Lnfvx+RvQXMTVpqc9
+q70ocPRp73DoENEkMKrBTEsztcs1lf97uy3JQVBJrrlzF9lWud9mofMmzXFFJAfiVC3FIewFOC/
L5wEzGcJ+VNnVjnOgj3Yfjc5JSrJyg60Qql/srNIVcAo7JtjHagKAZczDPH8VVkKp1nZuQcfUecA
aq11JD8uPGAXMBoFvZc5sIB0VyFfJ8qkI71Td7HNBHmnqKUveBrYKjIl+KBf2wiTBtgjCM0H8o+C
qAS9eCyAPaoh0SeUSXNGWhJxHF2TDz1IHTJ/PTRaG6loqDNnYHlfMgNiPjXuGYM43NmHllSyBj3W
tdUFm25x/2pxBO3Vi4GjsLG/nJtRH9BNyjbu1YpUI2nRlnsXZHUvG+I5t4WaF2Hc0kr6u27TmzJk
a81eAaJGaQ3VbPHG/QwzrhOUVgFF7X9ZC3uQ3oJQqrCV1YUFgsYwKb3BeK9quB40S6V5IOFbb0Yp
fvzAXwGk7N0dqnCdqobX+mCHq0sSJypd6kW/4PLg+wZnkpqJ2PU2PM6c/UWu252cotKbFMsRY3Io
4/7eVFA0Vyel0vwinKnkkAPkBv9OtCUr4bRNcgODgz6/rvNfg3P+L4xPlYzeJUc0PbnyEnW4/TIS
TnA+fkBh/U1OvMjMUt1/0ODueETcLRlwr++D5MjU1Dcx9x6e+wKx2DLRCOVyaE5IPhXAMO4jIM+d
jg0U+6KWHHT6f+NkDbCGgY6nj/wH7Zvb+gEISk8k7iouGkuPspSqjP+KdYxG9LV2TrqVr9Bqp8SW
Fnb+Ml+rQfmAoDye+/rRF39Dj5OSKZ63i/uhtuyVRG2Iwu6MPF4pGqaLbuQnxWwp3zgkiQzo8QCh
/yX3CMzcu8lsLSy39mnK1ugsR8U8/VgpB94o1lM2iQJKaQQD3RR6EDS447VVWS12omGiOhq6K6G8
oIxGKgey4tcR8dJhY3bRUVzo9Kyuqf/m2H2HeNevjPMTD8HXQzn1I5MP+1r/RH5eA5BeOSlgCZ5t
nbDp1j8NAm1pARguNQsSDgRvE42OG4qpJrkXyo2KJRT+yfvGlJJJ0rg77gspHn223H788I+tWV6b
141czHwXIqyuUlAFIePymCBBUDJYck3C7/bVFUOtUc1HG4kyeG9E0TbyIZF8GlRmGzifUyfEUY2+
RholrIUrmQYATPIhBtrOqdXXPL8nvPcYi5wqVFeOWeBgGWSIoESl4DqLEMfxNezFnAVvOaa441Fw
/dwW8BlZFJlIxJx6E9i68cuyNmr9iVQzL38d81L29uGOFabJ4fEXfDK2+EGzOnjF3Hx1OEt2IEuq
o+nt6+2FXjzwbk9xtqmdD0CUTagJaT/BNZrJOd13p3M2wi6d/tMC/kbKR62OkgglRTTWJndM/DnO
arGcDrA86qQQLXo5+9ZrGKe0V+qngVt9Xf/OMh+lYBJvoFwnpCY1l3EKI3VdFskhujQSJrcRmtJ9
0fO4lf6TY4QIdn0dBlxL3laysIcfK/srsVRg2X78SfC+gG/FcvG7gb59Kcx27GSryQ1g+mOR/rVa
sh0xhCYPT2O80C4/MtcjfRoR+EY2nrqgXDmGKlmT12PVlIbtRmJoxtc+RskGfwekIsntJSZ60LwU
kDDSr/X2R89A4oQq14cMqxvBKkm5szMr5lBza/xcSVtclrJKXh33t8EFZLeAxOBGFOw72zDMdU9T
NYDM1rSimNRsGyqkOPM0L1T+7TEUai/TDmzDBY71Jmi16QFqI0CG2qSwriRd0Zmp3HmyMVztqAOe
hZoKuYlQRepLItMlk1h3AMlxM4XZ9M/p4hPf0OfQ3UZU9QRSaBpWq/WAx4V2lIBHB/Z1ffByT4lD
yXK3LGeUeHXz59da+HGWmNLZOS7tjMZqQPPr6sNIEbj9/5AsaM9x1PRD0usybc7KuNX8RkC4y79k
L9DEXpcfBGCjW/cK/BWaUketIJQtgXY3bQSZyvHVy1gGMd7128IhODZChg7lLNlwGr1iHBxxw96q
bGeVueWW0cUjcF38OTkhS4D6b9SVacMVg6+hMsMcJ89CbskUQVQhyPBEDW9DH5wmk0XDgncVw7SQ
3yunJYz8ogRBFPcSNnes7SJBqV3xaqFEWZwsDSxVNdmwMxekowrNEzuC5fEDo1PFcPrOwfVg5DUX
uu+CUug3KWUB2nC/Y0tni2sG6KPUw+4q3Zsr5sseUu+FbOVnAKnAvD1DcYv8yC/+WC7a9HmcDQ2D
ToI72IKZZ72KHkgo76bsgt8HwvqwkUj8/RRHNPsalpAf/UHaI4hz51N4FIJD+HFNc+gdBMMhTSSV
pT9rpEpaLFm62QQQRJTxqQwE5B9OSV3y0KRoGnrQ0AXsErCVBV4JsWzXKxX5WeBL4XW/C+QryfHx
GygUloOYpZCcDl9mOAbIKRi0cy1NzmNhjl2dmtV+42+dX2BRccE+E2Vfr5SFHiKEJyr5UH4refE6
/NuSPXv66GLrEZPLCcg9390b2Q+GKX0P0wr6lunG6ijF1CIMRESpDr667rRLJ0a/SzuvlnDS9hKx
rVTtXd+gnhOGlY/wGvJog4FkmLTfwT5Yc95PdZzJ+t3swglC8OI8ygkMaRIkgFAHrY3WB4dsWcu8
QeTS/Onww3C9pQd5ezLx1TF/4bJiMi1TgkKR3nQ9Jg+oafI1CXu2pj1A7RJNP2by+/1xXvB7xCoV
6uNv9slCt/DL63b7e0XkiHWgY3eil4VEVdxz4Lws1u3Deqxr935Iqhmyk/RWrxIwE57xQwfkPChn
6AJBy9B20cJ7TfigKx62zsvtid/4ig9S5qkRhcTVvLeW5cWQIz7Pf02dX3mVmzQoff1Vr5u4CqqQ
QXLhD+luWbXrq/1DD9Xq81KiEBrEbsXb0iuCPVo+XUrvpl7sODSOHNMTuXFE/rHCKKWIAjnX9txj
qbis+m6iy72b7In+RgXW8vAVL89XB2H6k/n2VVS/uvIltZR06ID7RTbd0uukly233cZBaZ2y5zjG
hGJFvZdNNctpuF0GRHOdUVFkGDUI2aA59+1MNTIU8mU8YeaewgLwZfR6KXS/IBhSv0j75bjsm01u
RimjHspfScFFPBIX7upg3J4rLtucUVTU1+1m69mVTSzOkabgwW10YCumh/k7pKB8Q1CJQoCtX6lS
F2DqPKuifS+FTSq34t06kuhWEC8O7/CGWurA7k5RoEeTwYvoHG1006smgS21BY6ZoIVpEne6IyJq
hneoRwrjLrSrb20hQEPu6Gsh7q8jxx1D8h6CnqrMrYNz3u/W6FtEaB2u4Z+EA8XE1jRQf7wx+HXO
ocD62N/xIk+hxzhPnjrOpmJSGnO15FWaRA4gk9h0kLEj9JhMylJ4Id6GVHFvQlpxfqFWgF8w7Q4l
7vhTZYGLKyBrWxOBrz56TLlUrRLwb9MOp4k5lJeyo8a5yDqF+88GKaZrUplTZpWj5fhLS88izdWN
PcaK7y1LCf0vOq87gJ/RkgcruWBl0My00jigXcFC2Aw3d6vWca4Rv2llTUF5oSwWPwSUIs2qxUvX
fiBJ0gxdb3Ghp7mftcXU0ZtFvFFHFx/kN+r+4U92N8DOZzWbT0VwFZNmUY4Y02Jwx8IciefU4URK
A566zZLssrYYttt7N/hZEiAHvG+2trZwgM8diHh5NmFg0DYrtMoYgv74ALsprJ7SiWJYd+hh8Isd
kxcnLWQSpAGYagitdajtaDQiFYwHzgbGma4I0j6e/vOgUFnDk0LPAM8ekyMMlU0KnNkbPdw6aqxP
cg9yNg1XwUdrTSF4GhYB5z6dBx8oXA6M2r3xfGtevYd6Rwnzfe1NNzKAzxlftwO2qorNIiVQINRO
UuJvQL0XCGagDGDsxPKoVeyLE4f30kBkOK93CCg3u+WXaE/rWYOxovjmGN9mIfSCmM+zh0efpUEN
unc3LhkYAYBoC+fX3t3aAjPmETRL1uNavUgjRbAGjaQMDys09xawyQnEQt7OjdQFKKBb8pJtPgMz
fmTvqXZXWE+R5EVso1xlG9L1234IkKS36fu5lUAysuOG7313HM+FqVr1wCLKByc+hRTQqsLrpGmi
VQJRsPxRvsx64n3t4JcSvBg1vxjf81OgW8yVdevtsJhx5wBHU58udp1F24fl80MAUpyWTGb5faFd
d2fspr0gduVNMVOPCgLXcD39l3J8T4IoRhjQgrsWIq6dXAhbTptx5j1DmG+54kIhI3Qxd2J2YrX9
RyW6uuAmRhLoJsfnTeaKGLOi3wW1WSCbNkYivjHnabCRKWw4jynimE/SMXEtIeGkri5RQEsxIF7l
xJ7TSECYQNc5nm4IqdckA9XArd3wkFHVffKNkTmuYGUA9rlq8eBWsVfXlUEaks+KnCEqbFnr/abp
Bp6oh6JCwXN5/1RyN6ZaaIbQJUIgmy09smhV4uJGvlxns7P7oobh9TOzUuW2GhuRuDcN0eW5uwy/
MMLwnfdQrfvtgw6rnAUjJVN4NimRGDnJJzoBrE2dvdPYuC8WJBJYWUC/nhSXrMkp8Sem6O93bc8D
HKuK0Zg7jAJ6o4wKEf1qLSk4qQxGM5eu+cJugvrXPqu9aFRe7drcLjDoQLQKRiR3kgTxGzP+dvDs
FCVEqgDlsHDMngWgtWxE/9+KmtJBvWPNSRGsKMT1ciTCORA3DIBfVnSaOGyAo1t4GssanZNyh2qp
A5C5dPxgBnl6AmdlprdMaWdcXj9S1V0MAcXDCgxI44dEsthXIpn3bFOFBXTu7y2GBG2id2+C73fg
vZGR8I9dnq48A+fgxzvfTij6Ag5qie8x6+F4CUEkSJjnSEf+RdYVlOp+LrOXrxhqk7NRVbXvE7vD
q6H1jmX4s4x7cKguv8YWKiXL4jZ3DqbSVl7Wl5ftjnRDjK33xXGVcn858lkAJwJMXNFBWyLOUx4v
Z8TmQEJkZf9wslebgEg6oEdhgYFvYqjW5vi+sRFeP67cFakPH0A0i2PzXqBIgArMAPgGi+cL2D4Z
UYutGrcXo6Wg1fhZVt1xVOc4knsTgogdC/6pd8POBNHb0Qao1DS8gHZu5qlqUUXBgmgrRr/PX/h7
GtxWrVtST+gNnlIiOOXPR3WjCvxZcCfQdziCuRJ8sNseyUEE6BwyTjBVrLtNx2tSKImzdVU7Z502
nDOagyQFcijrm6TmS3JsZQxs6SJcPhWB7UzwejNno4suOT44w4iLq+SqpEaMXKdvnGT6XJYSWxoy
MRzpGfGvwzbMhGYfWYZ+MzxYErXQFzl+SpPCtEgCMd2Q84ZFQ2RrHvvIB+DemPeCziCJrlfJthwG
5YsSkUx6BkGfrQef4JgHvN+ujpZnxTbHvtGRbpB0kECveJIlz5qJ6+KnyeArUkqixp5WiJI3qV9C
JJbEi2s1ls6RwbRJNwVRq85eoibLPuSEuEXI/gjZ9cFm+wlwqeSyF4M0/CHyGtaDO0XpstxDFLZ1
FLJj/hwys0f+xaPBEzau0tyQqc0USAzpL2jMgfPf7wo5rVR9RheGBBFWTvqaz3DobZOt08ado9g8
r0Yfhwv4dEN/DyO1/GPzk0olwaPTow65RI3VMkeLsZgAplg2ay3VJa2bsaC5jsuKPzdQEIhZm67R
ds1Gt7t8pQxSPbPGRmC72GOgw7/PjGsX9UBM3ooIc188oVEVRca9TGpWq4DhZeeMERCIK3e4Oh/n
XdsGjZ/01R6kORjClQ3UO95MLieEDMn6b1ubKl0fhQDLAzz2KIuDRjddhVjRi6eK+15JDk03aNDc
GPJdUqmyF1Yb2oOCQ35sB0gpxDutYOrS5jjtne+wfEnFeBROkfNsHRw6dzN6EroBSr1sQEIzODjV
V+pfP5MiUR9Dp4dsIVGmWMtK9Geb6/HtSik2bHsQLOHnTo/4Q7vntxB/Po9s38XEzdBTjCqUSy5d
PRc0tX/cT3zU0IUucxsN7tDa9U0zeehgPQeIXlU4ZQ9E1qOehkZErGGLYLr3xcG3137EQUc4JFKk
2rWlKA7HD/qYzNJMHOq2eg6dliE4NzNMAksAP4FAe/fEm3jf1/gFmTAUv1nmk0eq04pmCQuTENMd
fqaxUPE7Qr84oSwTVCo6ZkO4wbdu2bMV5URpranzO130nEdyaX0TsKlj5hwEIet3GzFgau6i8I8y
n4smmTRYsCQrPcuQfYlhctFdwt88+xkGLq9UAr9yccLfV/K16YNNHdPYUqSSH5SqVvk5C5anGBXU
MW13PMldwMgGZOpUxEQ75jFY+UvyzXfXFzB90L811iZhwAP5eNJGyNEbfIjTyqbknMUZyK0pdbhZ
S93nD0cyJN/pfC/hUcjxJDb6871wkXRngWX55kifPeXIsQyddquopTgSmCdd/4GUPBoDD1tzEhgp
rATNAoewO9zg3Kq3zfFlHpBckecwls1L3FVXCMoYilBhIhnIKM+HYygogeicynHsrVfxD2gXr5xm
a/w/RxsCu1MguMtUj5nerTqbyyLafNOatzobUc0zC5tkteG1v9wS6fG4M4qWbviSRuRGfCNTYKrR
FK0tZA2bvaNpF2LirvsSKEL55wwD3hLeRrYjXcuWCD2DxL/1l1GUIf3yClyzWJjyKQ0KAvQwFvuL
yCF0l4o1GDRGjvZQ9DZGo6bU8On1umrepDKkhnkstECGwNnCz+d7S/v9IiIMyWMjJdOcQbUW013z
xqAdF5mrxKqxS6+YsUjFU3tPP9AtfsMGWFQUjdooprAagXgaaG0esIzCiYVprDD6BJtm4g+JX1ry
fFsMa/vfSVHxB9IVm0RjD4rg3MZ/EOu/+r+0DJ8KEa1uGPCksokC+SVNnaFVKcL2tQs9uzQdQq0I
CHzmYs1/4mMntc7bKUp+/FCIqWw7/RU3AUM6ctlIvCrdGRSSNzce+hSgmTDmBHPpk3Lzw5Tx5pUT
ro89IwQM0G3AQ43lRnVqKbjPxP+rlaTwzB51ov4fSAVX2U8ktoEYsIz1cXNuWM4gumyXg5pvSyb8
buAsXTTi5dM7bm4XLkOMWTV/KLTMdhUQVpFuP7kFQpUG/mIskOjPTh4a1HXbbEsZukj/Gz2nsKo1
P5K5Fje4jWrd+dkNGrKJ9bIlzcpRXyYKfMbJvCFOt/prJkiIiScHtlGqKKZHHw8dF8MnOwveOtc3
qVopbNQiOWr76QPvnQDGkE624j901YgRsu/aLaiuvMvVg9MM7VPvo3EbIvOA57PvfiYSPaYXA+2E
bJSd5p4ENi4FyLy3DdYpNaaiAULAbhkZcswdt7CfiJ6i5KMK2KGAxzfnDldy53fZ2vlGVgRi1B0r
swr+Esx64t1ndvvdOsznwKZXaSfUqf5QtEaZyads1rYwcmiwL0KAAOVWN/cbRUVswuUEBhNGt0M+
u8qJUiLv+puglQKv1CnkVwRHdNqIFHxTpc7ArK8Lj5FWr+c+ySKtIiRSTdHRVT5nW6pTUMJYeyEa
FuraTypChhc0Cy62K2DSSU+5XJebAtJmOM8in7PCQoEL4rKAnVRbYuDFaUiWgu/caQv/HmidB52R
OmqfbQUItfn3CgtUk9rFyUtsDIaCilCnswTwunGWWk9KJxsUOoINXRUDDc92u+Wh6D+XJX+etlOz
+eeaVFiAqIa5ypogvT3sLR3XVGZpRq5XrU15N5uaTokT9OL/bIvGIMz5GSdxC5gtKvv8L0LGHGOm
/7xaaBKW4gm1cQlD/beP8EXRtfbkfQBpkQQA8VfiXPcBt4mhEADomyVq7SDVcgfEp1gF48vAa8cr
GygA3uHPlPU9vYcFkAkLP8UZd+eKN9kRREJh0z6NlJej1eELi7URn+f6DW9EHs8Auiq2Hh2O1Qe8
W8ECap47TrpaC4s4Fu8zMFJ0nihNN3h/OV4VwxpOIzGeUV06suBPbX2SNW4J9fLJ/8PVewWT2s7I
6jAg6+55GJI0Lu1Cw0+J+Xe+ipxZQHCZDRhJh4XaEkQ7yBb9/x95R4brPJQ7K86DXttPZVkkAfym
0rgi0lPb+26Av0DynKwBV1uk7QgTUy3nk0ESJYSGnm70ftaHl6J997SJJov0VB8pujC9ft54gR8s
enYpClvqqIAad3sLZh5lD++jC2UsDi1LOWbrKLsD28ex8XsPWN5mCx0UqVvFc2cTW+pX1EowArXS
LcSAFSgCznpGf9RAERozciay2MGs6xpWkgvhb2lXir1swLIEz3mfirrFoavQ/g1iWl11nXGNW9dD
sJDdlOB86JXDegFn/WWWr4OSeLQC+Qbl5Xlvz4rdpYD9Ml6Fajd9ltcEbeGHyn5PuFaFLgP3qW7N
/t0nViS0B274C1g3ejtAPoBVEUzhrUKSaX/2VUGnkYJB9BlDXrzxTPGsoL32YTVvaD9fjh1f9HNY
UvIDdMdaQygQ3qj6NSuhvzdqdIWmQQMXD7oeubWqONNoxaW0+bAbO6fZWReIBubcGGq2Scgd8yep
QULCSwDbWEIcLbISUjcD59ZnijyYO3M+sPBf3YHOb3a6QSTJPa0fBo1Sl0Rf05VxZXjHxWykVHrf
ax6IyDVqmRZ6aS2g/rj/YniQGeoFMhSMLrJF1qRMWAYwdplpWksuka9Jn7hMOWBCgbuoImzkGH8S
3Quxdc9NRE+2uB6skbdPuu8V2pZejBval3vAeNqnahyVVDURufhFzlM34UFxue8VrMfkiE4CjOaP
aZYaZIEVuwm6kcwG4BSEOmJQrKflcJBhu/NZS317797ehyWdGZl8QDhvuIZuq0tB4U2GaZb3beZb
ib+gT7QYFEeF/hKMi1Ghaddi/kf+hP9gWIdMJCa0p5JNY2qEx3SArhKlDodO32RldQ21UEmMJrBk
aYBmTApZcY2N8NmfkUqnfaRLfkVT3MWvWqLQgSolpzSihsXqPWurRswb+NC07ggTPzC7jLlwT/8H
YBLo1NGH7oZuy+ezV5dV5JEaRtMhbkXD4l58rRAga1ntgK1a3XUe3bm/WdQH7M+Gq5OTaemH9czF
R86co9O5+4I5G0PaX8LKefsFDMd7ncYv6eY/QaN/B1zIBQeLCDef7YA0jMulnF/8LMGYPFZ8G0PD
echay+H1INXApnlOxMFuHaKw/i/ytN9wUpoF57B89OJBchgePkMaquLAP58/q6Nr+PQ+gwo6LxWC
BhxwTyrtSEX1plzmUi2hGGqx5/Urm0DxTClBmpTgMVWI5igscifWuHmi34UXR8WE4pwmaPhzQ6+N
mF9B2Io6McztuRpP4kJtkqQBgVDikRn3dvHuqabXQNdyDOMwovujPu4B9jkEtySVt10zQtUnB4xG
VhBPZHKcjjKRekIJ1TMILj67zyBdD3IRAXAOa9E9/Q9fa/wkCihi6EJKnhursB+SIQY8HrPQrGNp
bu5GPosU5QamEsdQj9FO28YZKvTpDsLeB0Bqh0q+/X8TJMWFJXuJ9LRUVGRfBWrJ5PIN0Shcqdrh
QxMW32ksfChaizra2ojfo1Jt9cpZATSDmz2j8xgWVDSzHtoQDD7WXq99SLShST7F7r/N0LFDAbHJ
KtG22oCVN/Wxt97A0aniOQ/pJdFal8WJy6bhOh4dSLMz/AJfmNRbnXulXlSJQVZWOZHSmPbCGeVz
QSVKin+iLzqlMga1nslkfE+WGkCLiCDwfEQoc2K6uoIanjQ0ZzXioixSTmlHSNCXLtj0XI0SCZJe
Y6N7sSdNB6/alNiVLK0+bs1dSan43gRtGgF9aZmyDylGGZ7TOzPGiPOqcC5uZNjvsTE02fLZ1aF2
DQ1gK3ksbYkUjoYrHHwxf2YxE9EzwKQZMmzW2Qx15jXjOVMeMsuuC8qX/E2IMcRp+bJT1P2TuwLX
jxeEXtCQXKApMiQbciGsTK51/w6VaoBAVzk4ZjCyhZBp5ocECAYix1s5apGTC9FzawTaObqxwXZe
Z1bn96ulN+pgMZQCSF5kX+NO9dCSFrkRGIo/UJgCYKGHuALkWSrNEBZ01d6FteludHErH/XLzKyS
wkJ5CUJ5QZZytyt7yt5gZELahZysloKm1gKybEzNMJfbciQaeoa9lH7z6hSsG/7IAE7rCv53DOYB
D4Q/NKRUwOyvwci/lU8kH/ZMsbB95ki7O9YpQDOPe/TCD5qtRdVsyRTXQNUEDeSRzg454of07wg/
K6YUJz0U74YM4Q3UYinWENos41O+rPUTYmg4y8V4k8upBIbXMflG557ZbnDbgX/pGS+dmV7ds4k6
IfR10ihgAUK9M+ZE+9iq28/6Q1hgqdXW6rrcMywkgujolYddrzFj+LZXSPWcR0LwWwlOV8O0VAxr
9OfKw/NdlGWVHzWphZHB6DtsHc3DPGreNhQA8RrC3qn7WyN3JFuamOg3VZWmyD9D0in1nLek/eJJ
90XVkoAqzbf3hIkxWejmIhqtyCtiB2Usbm2ky67CkNWsz1NbYJ6Odu9bKo6a/i05xFc3n/5jtx8f
qxp4/BeHW1ikN9Gp5zwtM9rCVXND7SrpxVeENC/AVV5jSk0x2QS7y1ojimCynTrW2KZRWR9kcwWk
LfTQGiHjQdgGG1UN9Cc1rOLqpUQLPMH/3gj/QS45ghruUuOW77gChlYn+Tffhhl2oh48lzHc3wah
iQfQY9QYQp6DZ7pqLnBAkqNYfjqOjc1oULfUe56CdTOW2I8TmH/9tOjx1qEWnkjdl9TjLF0kajnE
718fhWqWb/ohWFpr8zJkDzaHCFHRKg+vHEYRGTea1lGOYtp4Xoj9o2xeAXrAJMbPdJhHgk4PhRl7
FPt+4cQfvozF88GQG7CNTj8e0/NLfwXxkqN5PsmFITp27kJiRZFcANc8jYpIVIffSOeYWOC47rs1
KbGbkz7NRGijEnE7CB9VQbmT20qpPLXVztUgRwPmWt0pueFAyWZ/1vAfmxIrbSPGIYaCCbkBA5pp
iukvwEFXBWuXbMtzAg9nDlCPDWFr1PkmPy6q17qG3Q2Qxr3zyozgcCxKIM2qeRDoBNvOcq6SZb2b
mYJC53mAiGmTCUh2jJA/MHoziDO3LYAlHttDCrEHrDp6yJgM1W0fYuvil6DvJHa48xYFgJSBq1lN
Lzb6o/G9FczTNrtqc0jkNi0UUkkbicF9IuQB8IwQNAautDFCoOBQJrKRlOEr0oiyZV4ZY45pOVKt
mcM/nhbU2j/Te5FhnmYb/vZZ3eJ1sjvxnRvIBBMuiUHkbs4DGjQgOrKm/Q0Sa2dyQDIdPDToLeO1
FnpYre+9WFudNBQivXTXQXT7XpVsWEe10qJipa2XsOSFA+1C7ItRUCBY+uiXVlCiCwxMlAkcodj8
31aFO85/g2D1rNnTKWWMUG2UpxynZmg2HESFgG0MCCJ7ZE60DoAELYPLcKb2MICAMbMHgn9KHZ17
dQjRDJfvhIeV3X34E42rU1yxW7lyXnI1yI0BrGQGwTiNDiVpwQ/PfsX9ZycqO3KskUUmToas6N9/
hlAJjoS54bJTyfm3Ng5bGgbD/xW8GegQoKgVwZbS0RJOrD7DrqbpIQZQbRu3mCijjhwUZrJ+71bS
sumMBvt5KkHPvIDoqSMMua2ER29b2K90UBVuVHGYD/m34RkBXP7Qm38nlKB4gQDYBrHs5xACfZ4E
LuQQTpR9qXwqZ2rvp49gYH5Mc8O9W+bsUDDHvvGZiS34Tu1MnzWJlYKEc9QynbKeRvCvt2splzCz
V5iczuMfOBSqunhy7Kk/6u98ayVPmsLBRg0VgVn1pyttEWyIJu0EE7mUEYdDx+JztkAuFSCBHTYs
/dHRw8KPxS37HRvAW19ZQ9mqDforilaeq9jCbwj2tC6w4YRUtZ9SEiakGqqcgk/qaE0JxcRnjfh2
VlPdAjC6Sv8AIR3mMCpWK9oLRpw2ZaPQscve6lIOPngZNE+bKzdUY1jp155ymysClobfIzHBOItx
bds89HefrSR82W3g6RYLuc1q0SfXEKziUNvfHNMztvkB7czz3CTaclQ5uq2mdXdRvMSRPfduLIPp
01gZrO5yHXQ/SqLsrAz2HryDIMGHU5KIqd7sle/pNNzSHIub/dTYuckMJin0DMuahlwha/mHyCJc
GGV7HBl61okqikPCtgDWmyMpwyYNnrNyHQzOdL+T8ixNVvhdtXemBgcaK5mh0Gye7MLM0SBg1npX
lC+S4iqYCN3Y8fy7ObSW0teL2sb2pTvxB5ypgRuusRC2sx7AeVnhhZyxwuGxIJP+EfD9g5EIynCZ
v51fwMu2wXRzv2vFwc+WsmQqMMaSqUhd0E8q9qQ+WRP/b96Gy6HFP3bJJPbeK+K7YOlj6/yo4Na4
bUGpizT2hwrs3VUDhDa487yT9T4XFrXgAsoaQgu0cGpZqoLbKJ2y+2BXO4mBfeyqqqrJmP0ONpEf
KKaEYiwZgEM08ohsP6yPpkMWeU7TlWFfxvNa2YSTM9pUs7shwQ3OzPSWtDQp0pvfgHCVjNDe3Exc
pYdjuCfK9p1h4cS5kjvjtgMRj/leRyYAniKVXYFLJBnJ+7AGFNSrji0jLumOERhzPetuBnG6zMAg
Ut5eYAepl5QMx+iQ9Lb94JwOCd946O/swpBeLPlB1ZGTSa008A3oKmlng/r+4cG2m37j8IbeTl97
+pNs1sgK0NMnM3991BLbiPwuv/17SHqnbJXhtSnRQaXt1cHXstZg3nKs4QyKpYbueCIwCO/2RMce
Oj69xqISLN6UwJtHj02h5SDo318dhrT9lrQCt+fPIGfA/F/KYN9BeKJJ9C+VMbeX18MUuagi4D6p
RQmX+t3Y0FxqXTUBLy2/nmZRWiy7HrJSm3P/L3YMBz61VvhbUt2GV9QBppuGvT3rdloRnNIk3r3e
IvtSjp+oRjXNCRiKiMXMkT5kkrxADRkyZszzzfyN/VgAss4mtcxal89h6CnwQRWiqHhc0XS0rYnV
vhOmO+zO4R0w32OJJghujcNWk2HryeIEUvSz2DODcBa3xwAEMj7/riOShqpuZRbhAncPVy2IwZql
kPwH+wqJi7DySW7MMFOZGNaIrfLU6Jf8HeR3hE8FFNnZuoCmayf8hEWXH74PdBR74f9fVd8sk/zD
/o+GMF2sFer1sO8ZUDfBEFNDV1QRSD3IvA6cPVXh+ZdeUlvMOae5PzKS9edkjhD6OQqEqxeuC0kz
/7RbrSlHyV7QcEmn6EV2+nfaBA3WG0uT6iEPVunhZYJEQmS5O5PMHtNVCudLXEn5+nRmJ5qAVIqz
wgg8+eoTKkkwTQ2717n7v+ZzhgpgQtFKrWVhBAcXPLZLg/nK9pDDbwWvUupykaun5me3qe/8GL5B
KiH4s8SH6O9+ZzXA/KlIlxcsFybBm948DfI25Vvw8WC5GoAzyIkBo74tzn2eFfq7k03KUiUbVHW7
8901FgPDOpmsldDDQZneSiFbvYbnaW4ZefXc5AHChAFAYJt/XiDoxkb454/08vFOUJol5cHrOS9f
yYFigj2AHxPVvpGIkA28n2hD2bQXKNPNhlnk+w1vUR5eFSXvIN94eLmX1o3wvxtg3bBoMrlq9Yg7
r1pjzCxRpuBcI9GD8eMJuBel9aeXic6AALsW7WdO3DqElMIPw8qxbzcUiOq5Kds9lhznb9/xdG/q
+3QeohInEfGF41OjwQQidaxXnvdR2skhyPjzGw3j4UJLhDO2GYBGdiYWnSVXK5t0UxFnsYhSDYHd
gDJTa4f4Ud7Ndd8YGx/RnDg/7VnS17XFFJ4klLve72NbJlQE/poQ+F+vWPwro82JC3gT7j3pp4+X
cHOETtkL3XyTb97kSCLwRLwVVB1XUl4PvOb0SmGbt2lbyzzhmU5nnp+dGVGvTFQe7gAiBztb1E11
cLtaeDcuvQvUmXWQnpGu9EXP50Eu8n+mj/bNvAXmCluRHuXc5Wq1NXo1UEtQ4Ox2fQNEaH2EpMrR
EANGBTZ73i6ZR0xULuhbWpyWi0D5Wyi6twqUO2lTgIFlRa2tLFD6bvlixIKtePlHIcgyfDHr4pYk
gzbQmZ25ri07mo0O2N9RXeJXCYGVfEjgyXrFkH3B/tGwGyZ4N8vs7QaCIX80/tky/Cd4W4V3nUE1
ZBNynHayYCnKozGIVJhnRHx0O48sjo1UlWG2ftCFrd0Em/IhPnpJlYjTtGdtLfAzu8hMWcz+J3Pk
DHARhkywPjKVGgkCtnLfuvIB0C7Ce1ibefkSK1HACIbzJzyQLN422tGZ/32FvYD52w9rKdB3J1Ms
qKEm7vRaYGLLPEEvwn+LKs0A3oVYBb5EzszhNGj9y9X/+/Z+TYwstRN2aqmdJDr7bXJoz5Bartlj
3NqajqrTO7MqWRF1W6nF/MKd4xVWmhsHn+mFXoYuqIouiEe0i88I8et3tKCQomwWH/2f4Dtjq6/5
k0Q5438KiYDkrGXdlk5xNUlRgMPOkeZHTk8KC48jacP//haNm4qYq94GwXniUlcKlwRcWLDIMcuP
rXZpqiz5dvrI0taKnuAiDsQjD+k9384XAsop2vIwJuQif0CseflwJN+qx7ukcoEHbPL9hq2bgaZe
OdD5HYT8L+JSj+91p0P7mweEY44fk970sBw8Zob2NkomNqti3SCTqYtu94JW23oc3kuVfO9wroXc
GAhSLn389udZmI+BAWG+PnlQ7ygb5HcIEpNiVNyWK7zMqSVsbWhOiHmTMF2cUcqYmP3fGYvEvvpX
1W1dE5M2YC6n8YRiyzWbuq7Kj8B2buT2JtHSdcNw47Lm171lFQQWS6KfCIc5d+p3T1g26W8bfLMP
rVg2QxLqOQ1SDj/KwjgswkkEqXnWzkzsNdrIXaWHMuPV+5q6XD2/16M/o07JC+Di2acWFRR9HuC8
Hg2hB+TAeFjKYiDjcrxJyjAwvDRl8TwAoZoz41zkupSGQfeeL1qL3NbxjjOeQrq9G3eo6fvfIXf8
7StD26zNiat9saL58ui7ciuZo79vSbjpg+K7B/a+4f4pQ3Ld1eFwZPfKoI3gjM2NeNgZ6EawcpLS
lwE+1xyxNDgYNqzAgM5SSCkLNx6CAomyWleyxGpsPeVq4V8VcysFzye88G9C/zptB8GOlPzcI6Mz
Ot1NYqz6EqUHv1jsMcFyjrxtDlICgnABDup/gv3r2ZJwmksX5xOIWCyChRH4ZM2pzzMkBXmDgFUY
NnZEC+NoFB/hcI4zFG5VsE5MSmRbqOcMmdAm3fbUtCFyc613lU+e89rfHibkL51ntj7WorGdH0hB
ZE9ecxja3LAQ54gCvZlal0pgxPKP4Xzy9PgP/Ft8g77Gx3WwRNzu7eGDQUN5j2jKuZlpT3qgsXjD
BqD5/d4Iahg7UHqKdklS0gTOl93J3GoklBcpdmNVMOlDbx4KDcG11CjoVl3GqjFRbEHXZv6QDQlf
FjcyOtTcIf1uamiOZ2q09AD4NtLltq8PdoihPox6K+Qam19oML0gScRf2POc5AoAgFRsntOcO0Sr
RF5RZRTab82YlH6pwrNb936qSg2Hbsm3JclgylPKf3n5hwdZDSL5yLxIT1D6JFVX1ZPSIotZKh24
cJUx5bUI++dao6L+Hi/xuo/MHtVWr0ctgKKka5GO4weLnwLADwrruBiGnQAkH1Mt0MND2jPwsqd1
kDw8vpNO7NevNJ8AKiXq3NWqg2gegNriP5aC8xI4igQTpeAmAWJLFtN57LVqF8H2Y4FAAfhGZHNI
5zeFTVYWVuSQpxinGp8wWgTMNoS0tIpQrW6MmP+7tTYTZvS14bHAcHm2QRRS4cOEQa1ZVnRpmWih
VbcVMjtYFNvOfGHNAhmf7PRWiK2/h6Go6t9JSI1M0KgEH4WOtMvW40V4lso2nsk0PhOvHhTkqKAI
9K5tc1bUc8JbGRRA9r9LHJ3Wo0vzZ0cDyZe6bd7ZaJysWZqXKWh5E8O6x+hd8Mj3McMwXNgbhzUu
aMp3cLrv3CZznHAqsx5k3Y9qIodUEy1u/UERJkS+xtjj5ne/x5SHzmER2xFyJasiXqRx0UQ/IPW1
ExsK5zimWsaTtrp8lJxqrrvGUYmVYExtftz2c4PJnAOGARWEi0pmcRaol+++q2xhdvjpKzZ3CqQz
Ct4/wSRRBqDCA5X7gfNLtQEb6Ylm+uyVECVZE5WWeQ31fh273db80F09lHCLIqNuheNhVIOf+qLx
TYDz/u+sP4GVb1h9mHbT7VrjqA9toHD9OvqwiI8UGSwgifgfOxS3ddlpRSNVtE+i/edV5IKRHF26
FJSBG/aYoeK/HlMeGDLrP3N+Y1xIxPtn/JxnwHdbfaIsTJn2aZ9RElh2VLhdHOovhZpZrXaJcJ1j
CTkQZlyg3phGRX1AhdIBNd/P6TyqyixYuWy0ocQz92ExOdXcRNdLB1WBBT2GDJhVz4U7xvYVs886
/lK3bUBW9pKFPXE2nUrUQcQlgHKlMkI5FOWSNRU3pTkn4JBUWsAfVtxW+cgil41Tog+f119YqD+M
MZMUlmLm9iLt34BhSsO9I9a7i5My9Ryg2Q5R57EfD7kei5Bozg/INecBI8/2Rba9P7dZezLNzd2H
d/VAsf61BT6ES/ekcMxyKRO5DQWSz9h9Q35kMF66lpPo9aygw1oAQFAS4jvnYxEIOqmu1Z5qbxmt
cA74Ez1lYKTMQbmxKu+iCCxLwBtOzEaWJKUkPi7dHDqLJCz18tpNDABzVO1pE/cqvXUdGS8j4OuT
UrB/iMgqs5Hz9exUm+zhfp271KDxhczkOxtOhTqb0tueQHq3G4zkTm4SmCdR995XEsslrXr03Hir
9asV/MmfZSyRQhoEqhjzOh7Cdy3cNg8WZJz7HWtX0+4LOzEjkPVeMO/BHhvKiwxWWC5kxnLdu8sw
kN7MvsWzeSoD96e+z191BrH67VdVdpJ595Vd+Xs2/wXWE6Zd2USO3/nsy8ZhpqmuKbZzJKWUEAaX
quxfSQi94mtQXJjUz09CqtJTsFFaZkZLXgpAgF4dPHvjUyFAsV62Om8Fj/lPY1V1k5hpanPv3qi3
Np6YJCzT8axainVAtc6ZijZGCdxjZkG274si4FuEZWOH5WAmpQYpG4oWqkfrnbaQnpnnBekVGM3T
HrLFLg1Og7+2EeCLhllAw3Ma6p8cq5Tv+l2WTKFFN/8wESAEUxCqHGLFgG1H1ppzx0rvIQn0pTYy
DCR6HlrvCTf2AEoBvx6/bCQJUsulFq5qPHSaKBaheishgb5AGbtKlc5IURGk/7WLQF5/4j9Erqbx
VIwekW1nTFuSv9I94+9UWvMdZblCSXY7QmGjWrqNR4uEnIglGcq0JeMQQYUmxUDJFaQYQ8tI1uAE
Yg7lNbGTtDCeciYrqUjTmi5kQsOG6w+4Lj0RPZ//vYmLlTVpoz6a9o38rNaKbBNG9GUbPwSJGtkx
lMxxxP4lXiPPT/59F9WyCBUNgonD3Yrbn5WkKPwGejYta/+cjETv9zTs/1AAJmeXbq7HXWXubug7
rQMYv3eLdJNj76rXCYM0jso/HE8g1MHcyvyd4h4GMFUdpd3T6FgXF4gRfMDNN2Tsco/yjQMJ/Zu6
rGOAb3QthEa3aV+cSA3cl48rDuqTX9OfTZ/6x9UeFclZNBzrpbV96SHlw+5kNgZRSshMjQnCHjBq
sHodMytAI/qxUimgrvDwKOxcGygyBEo5uW1dG6LwygUdE4e9Lpgol++NxiaLjtxBgfGHyvztdk1P
E/fkQttK/2OEzBrqWwYYqmxEOJURAibllb0OZKI7OZAv/S/hZSOWm06/DakQP4iP11VBjEiTWiE5
WxkwYLodituJ6XN0271KHArYj/IeW+yphnszz8N4z2OQ7qYkDEAJH2S+IlT79uN9kd2epbdxTk2O
xrrz7vvqD6YOI6u/CGoTUob7kLwozjHofs2xeeRm//9yPwalNXCsrNBxH7Wtm8msy+aW8OSfhIg0
TEIBsMz04WunCXGCILys3m4+6KMRjLnRhfF0JE0HHpc4irh4VMActy53c9KAqM9JKNk6bSn7VEIJ
bPatPapQn8Fq5O+JDstayUJMEJkIihbGIEhAUyVugEssQwi6u8zaHtWPUjOKWVqHaA52eGLKyo5H
INMaNhlhF5vOJLB7DMUkX7JOIqNIfJhmDOZhTqL2feTxC+5FnLRLOg3Vton9BmlVO10Olbw0E5dI
lfPizjXnaX30vIc23m0PYzFuhHDFVi781MEvA4FVZTbYLiFDs0YXfttMO50zMORvjckHzzV24syq
fquG9qYW8h2BCaT4pVXL/y3v54bG2m9rFXZcf64dsgyiTrOtchDtmQKW5D0qQ1dKDQt8F4c+ucUG
E6t1A8xZICHInb7Wzc+itOeGnONZKmQ3QhhDfjQ0nN1kWYXJ8dpGLhyBYsQOnEaxScYZcMregaKd
Kn+Ecg3FQn2onO9J/hbv1j8JWOZ1pkQERwWpBr06VUE/vT+T/wAoaW9XDT/YyA3F5+bDjxGUm2PN
oM8a6Ip3hPcRHeQ7MppqeJAekuDiuzL3GcXM6Y8la0PXYXMwrFJdwVyjxbaIR/9RAapl8WODffiZ
r3Dq+8Bu4YX4ojbNTSo0TlXPYdhJTsNJkYtUW3hBxgJYKaB8/FeDdwd8hlkrDcZLLqOtcS1nEdAe
Ah48rEtqCy7N/HjR3yoKLrR0qO1xw4gk3hQhomhts9mTXAV4v79uVerUdG2gyLiLXrDjNFklO0FY
0OuRDjSAZ6XmZ0PCOQcaiqSiK95dmF0Kt+b5bgrMQtpIu9GLcVd41teaCu7+aJnl8fefUCkNdhKq
zC7WHhCSIvuhzcXSolT5HH6DHQ5Yrjpd63ICzd0+MS3sY7goERZvddbKzZjkT0VFu5bnAA0Eq6XV
fzrJRCBTHXFIqlnTavA8ySsqq5uU/OhHba7EnxXZNnm6OZNJdBw0ah0XDUCLZeGR4i57eqgGby/s
yyEvg0U3qlByH+DJIny6hBVyQ6KX5oHzzSNkhN2BV07kAclI6K0+HO82qFS+WRrDgtHr3qto1Tsv
fNLPA7lVwWqyTSY/43TdNas0IzB3gvzlvXTA4PYs7Ug+4LGXJDtStpGPE7AoEwq5AJz2Dd8mox0P
8tHbkj9nOoSgcfyxZS+qAPowTfM1usxUKa6EjrXpfJARrUOp/P0btP1XU6Uqtyeps63p0WQJmsXo
EqrT3uZwtCdVYvkvkhxHjrYIYBcitwcgtPthkovW9Uv9IkHa2e4AnvJ38ydzsFDD8ROWvIL5CYYz
iOCFzMWfRnWfu1X0Zyur18bLLrzP1mgNNBDvAsV5E0XmazCmXmOnQrk22WnV1VAgBvTwUWVc+/iM
jbz9ZGT5qRsC3arwjQv0hxow9K+nuTgyUfFKTkKHwuvt6sa71anHwLv5GVff052aB8/zEQxQfxrv
U2bQgAWnf8gd8php6sC9C3I/Oo+aTj7XEmoanfGclwjBf6PwHrdOzyLdIvIFs6b/2iv80WW1VNN2
Jo4Q8bYW2fte65O3v4jwMFqV7c64Q6J4cL+qMAmwLEdQ/wtJEy78UxhozQ9V61OOG5joxQHHBtKo
0B9RonEHW+wciBK1TzDScVi2em95o41cc3Q/HSOKKuMT9p1H0TTih1nRq8iI6qwpyuAhCelT4q/3
iqiyiuE7KSG/Wh7nfnmp5R8IuknrmB1wXIh6Q//6Xz+WtY0IPfT+LW2JYie2bIbhivr1IW/aJK4v
aCoysoJutHk2VImpv24LFUv07FfR29rtg9T8Xt/lcJCv/4hu3OE+0/UmJJ25HwED5V5YOYNLwg7q
GLSA2SQ1GLZPRoi1LuzgrGGJGN9w8EIfVxb4SPgRO7tm3dX1DhyXO/umJhGY5eeBrjQApzT3JlLV
KQeO/s5wK6vQTA/9xYSnZZdsDql7jeZU9JHneO5CseNrw8ThcJRapKnIdOQOCnYF/1QfsV+9c2X+
KUg/AbJ976AXu+6NFOGFFf82cispvh/ZTwW9QyFO5Kya3SnlmjaXgUfM8IbH/0voop76AiEdmM99
2FckFh+c4UhTNf21Mtl/DwM/Sn/olyzEm6+3IKHc8C9UKnCgaYIQB/2iKg3reosqWAZNYPsPFycY
dGtaIHpF2AiBx/DL/gEXvLnW3THBpf3sjuDn2s52axpSF95DxkQEKmNe23pDb7MGph9bvN7e/HpS
wBG057YlY5oGsESsy4d89sINUdNyUOjqsu6zGyjC78RWjjypn5CIG7u7MHk7x9jA/RzYFvjDpp48
dQ26RoZWROwZxL8Doim89ws/JgSmM1uoJUB4pZZHLmnbY4rMhmdlGw0gilyRL0dKb9K25uVtmPHU
pDmj6etml5cSijhoPmh1Jz8sf9XGLMAbSg8cU3oFtSM7cScYCBx63gO07uVjJKZEmLjIXMt2vfWN
4L26fhJVBeC3XP57hsRXtEFY75+ul5U7jjQjnWlEpxyrijkLOnZmeOBsygjWluJkgF9GyHCm2d8x
B5GUDNuNK6umU8J2VqnytbWz/MVX2ePetjeymtv5R8Dg7Uyl/csahWbpuevJnWIlUPSqcllqe73G
7yFj7nN635E5/rrgubia4bZTg4x5Uq2J8eoQ/iwokYNBDLpOR2Cz44utTvOuN4FlAzvBQuMANmp+
NG/HGT/r45yXY5EBJbD8CVKHJPOyqleJhPSLg9prHX5UwMYnXxTXC43h4kIfqxPLjjtW8Ytra4Tr
8gkhIGAejH9ALfM93PkQEQgwZC/TGG5jD0VkPklIxvfd/lQFLN/2XsaYi9qYYBIuv/K5GuP6yT7Y
qfDbbi5dTPjwi36ZT0JUBFssFyKLu7IeQKzvf48tTUTK4eyaY8Xrjo1GAOEXEkFFHlVDSMivgepl
56An3GNErUSoAouZBKnkfm9v6qHNUcf6zEnxvyoBAmtbzksqP6FmTs1yrNhvwgmSZBRJOqrKlUga
n5WjzW/R2kcs7Cb6/ZcqrDUqGxyg0+3chkf6MW30p2oeUVwseX6JnGt166dq59LWihujh4AwxfBM
TcYKCu773+alyWy9vYRFYvUWKN+Not0/x3/2i3A3Wf4ZcCRveOS35caMfi1y8vdKEz3pr2S3UQqr
Yl2U3qC560Ptcm3B36MMBZywVhcTe2RY3ic3AF7hKLsgDrzfyxa+gAjTAso4WUQXTkIXnLC8o1lO
UlFbZfsnhgfr/4PpXhb9a/qOYPbZq039Nx1lXNKEbxkzQuYue/RBw4unUAgi3Wq7nONMqWrV0n9l
TQsTOkkNrmtfyE+OcK4bZ5itUjKfB1ohp724zAdNdUL4crICZI9+EI3yQhlfhXHAP6WVk1WzKB/l
oYKud/4p57kiE/W0h+M2WHUegmF3px9Vu2W2XccRTamUZI6etAadcWYAxVLkCncB8OC5mB6hZQwM
Vk5dLTf0+lfBuCAoMmBkzbAwEkaG06jNS+D1PiWzm4kacZCjiUcXkUm/ydhTgjYbkdobmN1rRUfK
Gs39KKOt9zSJDXR8REPPsXKVkAN9nJdTdDp3gSh3dDM/Falc8CLWsoNj/KUk1tmUYnBnKonl7vNA
UC2ZucURT01zn9+2YvpT0VdFByUjJNnyQbxrWOjIX77etuBqx8K+ogGQTW/fBsrSqCvtzE8dtW9W
NG3Md3SUkps5yxIs8YWE+JklYD9MU5xZ4f1LBCyxtNnhirFK5E76VnO84B9mBfNIE8D64HGxqUwU
OzyadcR2s7/uB9EYk5OcAnViFUo5LwDJSl0JBQlSY8KpaPmbQipN41EK+a/jhou9y5W9VYYJDh+z
SWAfY9LSNcGs3ZqOEK+JfCq/dkS0XJJfNifFqgWCsJS05VwfMlt29Z8OcwD2EW1MrLbPi4/XaPuK
lXTIgqZeEDNTwALBuaG6xRS62v21i77vFvR9yczm15EZf4nVH3j5UTUAArEqftIA8jUAQu5LSO54
gQJ52nhhsQkHuTEUD9QK4WRLJN3EyAr9ijL7914uWsTm1DZo/r4EZTrnEM3kmf677UxuJCb8aXSL
YLMG1o65MOwiFYkd6NTgTi5PrTWEwRwdXgF0qNKrp5oScpLfuKpBDebqYE+BZ3LZTTyE+nz51oQN
RoOOY47+Uvea/QMmTcpoEXwoTfABEChQk4fBagbejtXFNCdLb16TPu1vOTG5arqQu/S1hjRe3bbe
uICyF0iPtI2r4VFx6DVRCfDvyiKyJWpr8ksM81oqjwz77IYokutqlTOq2exYIbzyRmWKd7q0MWIV
tADg9+EOQpvjWlYWHIGYsMQeSgfCV6lhK8Iurq4DY+oUM03RyOLxSwMrYhNteD6pZO5Gk1xST02i
6w91zOd711FhQNMZ1HXt0xV2AObCAePDVkXUtDjre3cF7wOmttI6K+PBH93vz/EW/KWtE6vkLocg
VhmF3oTlWcMgvzCv2jOKAGDh4uNcti546usjkPQ0ywGVcB5A58EKJWG5JQQvSZ1al+dHs86XGZqB
cOlJ0WDFleEHH/aeA4QYRRs6w7X0gtQQJjju33P3EEGgKozd7/ryJDc6fFXNkW0Q9/zZeRS1MU1C
81Ovezl8H1IhmZEXga925KVrob+Um+ckFs87gJYGzSkoBO8QQeHI35QdmMpG/tZ6aoBiZfXrWWYJ
mfAqkMa51U+EffrH4aaA6i4sAoyvOasq4kFEhAtMriFV8R+ft6VFk3moIn87I/DXSCDr6ehLlILn
trflnta9MxKfQGjNfvspepgt8cGogC/+HHN6fV1lPjMwM+3MeRmP8O46AmIwqrRrei8C6KVl0Dhi
sMQdxO7Qls/h4+VbBeAFp3ey4TIuwc+RjGTPTkHv9Mh0FUSkARoXuKLUBI9+2HD5Up53skBqWPwA
MV8nGEA8r6N/NJgaaEWJCpF2v8SKla8Gqxp6KpUMA6rkiEogJkOmbaVD5C/C4eDJ2KMy4VqCRvSe
iHCzPBGqASfaMWY/M891lAcktzVAkNiyK8GUBDO33xtgqx+Evsha/qfTV22uwE9hqGc7xzf2ScfR
tPtuMkvQ8BOzsdI2YHUj/FfVivV0sHxyy8MjkJyM8MFE5aM4eR00lB6wtkzryzzspCSdw9er+v3o
BHnmbWWeaALWa9amI/7MxJhUZNt/AqGMAWC/DEwqG00pARinsdvzvrDtwC7i1BMTHbyOy1EUB56V
k7w/nR7OfwY7//0X9u2GnR7yCejF0v72aYGV/p0p13i9FvlzAiT3QAK/wkO8kr1Dukj1rRHvZ8AJ
0BnmtFp5FnV5Mi1R5bby/N3AcsLQk5rSE8XWrji4mbDuwwNkkLp1Myr+geWLvS9abRJFA68wrqNf
KGa0qO6BLieAkxImoHoIVOGeyYO0IKlgWzhy6bam330IR+bcZ803ukYA4jQJ+NrF2UKyU7gRMj5p
8CMkw0KfrK8Y2S++qy5ldahux20L85ieZVOmJ0WOYSUpbdRpEh/54zymjj8Kvsl6O3BDGz7e9hqW
jPB+3pJZlnkc3uCvPu85JhC4SYgOCKaGZt9E8q6a597QeidOdAyf19W6Y0O8IXpIMC2sYPBICtyz
vB65C13mfc5f8KSRvjVP4X7RUYYXSmVK1U08eM9W/QgPdUlsypv8QaVGrKAujXsLc8U3skQg1HvS
RN0jFjhmmVTy49fHzDRjgDVQ5Bxqhbn5hgf4XQd5zbEsoN8daAbsNBIHWONW615EiGHYMBBJbkK8
JAkTvq7ilzVJYvYi7OFFQBD5YfaxcWdGn7Th5RsYjc/E82udBGmTpHJrhoV12gM+0+A4bdryxeQG
W1twuS51Q5HEdjRZD5+OllW8M2F8zyMy6y03F5+qjBgOgOOZzhOU9r0WWEiFlZLzETydfdjAIJM4
98mA4Uy4Bz8nktlYJzBKk7LxQymn2hrDxFBed28ycAlLM1yYWB1hX43GBQK/8Jdh/N4Jj7q1GrME
HrIZ1CfAY58Vr1Y4ziysuluLgDpx3iQb04MDd/rUfqHU9hUQcXB54OPmH/v1w6zVP5jTQGoIBDCo
kxqWju9M+qNvjEZFJ74S8/IDd2jelKcFQSmWcI7g5Me6ZA3XdaVdqX+zYjekuX0WV9S/UJ7o+FaJ
/u5F3wWYFzXwrGjAQeOaS96T8lyg9odsVDkRr54FOkINyjCaCgGZNLlFQHkdTRAeQtnllcuok1oJ
1jUQPiQ+p5qcFWUcxD69a0vC/h2gYpMpOQkHROoYCCdgN5C8XAxuPaJro57ZpBoInIxsD2tdp2Lh
YJ77ZKjCLBmrv5umLrEswcTWncyeJNQSuJUN5J3A11eLZBAnwXAmoaaqTmKIx7QImHv5a3FHOZ33
5Cm3uuIRBBC3iTIA1gOL0Lc5AU+pBTANDVHnNMjF0QfFTq1A/gn9Ir+9g184NSPjguZjWAbMjXZ5
Y+gnq4+nKP/fYpc3G0Si7cafDlLIhM30ErWKML9R6xfQC+J+1WBTTsNpTxgU/BBAma42wMb1O4oo
EylTBueo7Tg0565vsPEqt62sIudErUF9WncRjUDcgGnh+QalQqEK0joVvb1yTQUMqDPlcEvKsnfJ
HeaH6udprVOkFgI83vPenv/kvukc+RyqnLPlIch2/h8ofWNc03KdqT/hwVhW0JAQLlA8aB1Ri0H/
V1vJe0D+/zI2UhNMXMKprMx3H3RXEVk7xbT05Kkf7kdOvH6t9gNHvVDP4ddr3m8Tbge+vXWpGDnj
YA0S28w312vC7zC1CUmykynW5AnYSiEhrb3vDNl8Zxa14MnNau3pSolhfd4INsNkobPck0YaGf98
qU6vFrZm4RS/Km325HIQGX0g7jAHyFRMYuc6X8loWBtG8+os0lqomI+08+6ueESLBS1WCoJgcWHR
AAGFPesnxl9yORBh6ZWQuOiLIt5Ir58pqTFS228idGtm8XLYoFUILTi6RuCMcwSGakBsy45gk4or
72rfD/V4dAIJPS5Yia6aOLedvTo6L4YKzPWKvwoxM7eZi9/TwTe9sq72UzmTXk/bP1zCc2h77jkI
Fnq3JFj9Au+bEr21m3KpzMENjl67576GDJ+2LsJ/7QDOySbBcMmC1jB5bdyMCWdIzpCb3kLOF1t3
S84l3QEWKoIvy15uP7wCLNdKa4rxAGX8fHOEZ7y5gTOtPvNQ1xBsU8hxqUMOTmQDr3Bvqk8U8+/Y
CLvyCW4UlLle050xZF1xHFe4rXpp6totTbgzMPXqFvwQrzUWuxTPgClIWKepaezEdc7Gtn9fDplL
oTmClvlSRB+VNeAhHK94q90iUmWZyGpjQd88DtnUdZT0Qwl//VKW342YMnwkT7NdF18GvLFy/IaI
KUtGNlgeOa4WuRNQfSuLACfC8DjiO/jqTkcU2RYFmyft6pGgy9tUHaGX1Z6oNde1w+OhGD/ce6CE
hCFYtMgBrTbxjjcHHhq5FNWu8kwwzOOstI8QiZCah2TnPrX90u79mjDJb4ryppNUETvw4kOeCoFi
RBHwtJbsLNrqHDn/M9wxWTUmwaH4+ow4lQtHE/UNLe5k9yk8dhGe3/Cd9rXlEAZGzVYcVd3RIr4q
hAUMpwpmfhyEb82H6YyPufYTwLnAXVd/G/AxnOgKOgJowsLPV29Y12vypKgzVG7M515WLjvqjSeA
nL6fbVHThBVauuJwL07KrpZu+SMMAPlJ3+flj4TD9xY0FF5svWXymjoNzKmr2YniYtuZPH87RT68
bjoS1XovKJJZm29OjzwN+jSKNU9uBxWw7pWVaAmYaVm7jvsplM4kizWrAf1ueCYk24Daba4yd5cu
h/6tnL6JfYz5OWYuUAOGP636/UlXigX8K1hZGcNSih6P1FNLRRmMDIqJ02oluwVdULs/mped/Iz+
1G6aFq/mD2Sj8D0gGRRPtU4XYhAqYMWperfHVhm13Rl/chb8PYsyCX7lrJhLqFkcyOW4jganNRkc
fpreSySXbOsGyAcRJm3NVmpQ2DSiMDW9Biv171FYqqFMj/NBwuaY86jkARL/p6uFkr6ZP6e+TQDY
pjdmo82GvUGnZvQXTWAtdsdXpfeKkbc6uf4fsiMcv3CtGqimFKoUhVcM6Kr7v0DFqGnmkHjbf3zv
uMTQtUaopJOnvLxhcnTUzFOlvgpyVoro42BdV0l/pzLlcvd9IQLTf+wCMQ6ZQkreD6CFzReQOfE3
cIQsNuUucI3l0OjwTnKfN22cGacPKWTuAk5H9U2gIE53irD9Xmy5nIKN532Ev2WvDQf2u84yXBvd
ii9JDflquW2pFEvqP0hqa2s1WUpkE4NCCBOHu4NTSodNaietObn63Y2D+D4TSKHDxC6CFsYKdUY/
q+FT34rNuJtITApZOzJy3zj6O4Qb500J0RhrKCKHMffk0waRSY7cLPdvX8AFbxN095H5bt8vDreF
AmJYHi2FnKEWdItwmIEjnQhoIcDgJ94NlXIQ30iV/1C7HtzSxqiPcpSgWAkNGoTt7JhBiH/futaT
pK97tMvYjeH96nZUD8YF1tLKT7X2muZQoKI6FG+ok4LgznFdXcz2wRmv7pfbUzNERxExpahzzwA6
1lSn1oadOeA3+3VpMG3oXE+t7u8iQG0VwAB7TEQBwrqCmdsSAwD4FAfTUzRySdOmPGmJIbJrA29I
t5ZOYtNgKxFYzckWE3+9bOvM7b3xpefsUrgCeEP95W0RNusHPKGzPPCajYih03V68zRbJUz2tHXo
KBjt1bQRPOs0XFX5gjEHDxpe9sYo86ILA6ggR5rmnCjvuZyOZrRci/ISgovEtJrphatLp0E4yb1b
rXzXPO5R3b70No63EYQawvnX5SZTXWuyrC5+BJLJ2Z3lHWYyHAS4dT36Y3iI+Nw553/Eq313O5v+
Q/EHgfZxSLtG3h4L7S/pbrIUVTiciit0ReTob6MHK4mZH+cLhgxarjV30EEjZ+uD+TKrRuph68Ws
NkJPa3NhUqX2jpptu2XStGQ+w6pvkkV6mi5mlgWjj1C3xw7sdYfxsGJw6K2t0zL9LaWkNxNO9Y2H
p1zSATwzKd1+4VRJUG0c5SHptDK+PRr5QLpA8H95yeIz5LRQNVl7307/hGOUUHDbM0bOeL1I1UZF
q+NXKr5I2Se5Oze6CV+AXAT4OqPJCgr6riHhVCUKZeLcV+2fPnIzk3YIzMH4X9dSRrkv4XjUkF2t
wcobUfSuaCoQfma75Bl1U4VKV/hMmO6f8UprLOJ46+HcgOBlwIoagHU5eDU0WpBMMcO3cH7zIMd4
lM2DJhXzkNvwqcfd9TtR20n1RGbImKvnFxtwWGhsAhG43dfkQlPkG5WXxGKBppPuFf8+wNHaaEqm
JdrFL0RhjI9aVC7QLPtWlSY3s5b1yJOYV7h3sGdOzf/JwSuSi/u8e4b1HvEg0RydpEIQj1wlFGwg
KqNFVP1RWe+4yS2ZUzuNwWF+OgKxEsVTgihZFmup//I5/hvIYTDPsxO9SN5DGyTbCD7VQ5Pe+rZG
GUPvxNaKtdlxsu2nTN1UcZrUQO9n1cdnXtXVtEoJZR4fOOobWQZZYFBn2WsIc6ogNX1D3OwURzyk
fCrRs6tbKKuTgLnjWnjxfoJYlNWg+2zVsCtDEHesvloXARWQRSGS7Xk8ZPb1ynUQsH2S7enlpHDX
2miRZHhJhML4+iLMveDwY/88E5KvCYKNnd8ad2NyKavgnt5sgqllOmIHVztF08FUdF7P2xfemXw2
Vm7ODw1iWzUqy3qrvYHVOq0rZiV9M6ePAGi/L+1vRxfMQs3syr4pkIrNpgx39Wdjx6CWuoHLkHlF
ek3SHfc3k+JEpIV4NVV90g1aDTrjVU7oxrs1Lt6Fhk0pfyUHCiHX2rjTlGStfl2cQ1lbbCfC13Yc
dRHwBN1MXbhPbo/OJ067a/tqMnZbftJ9/jfFadzk4JaFNlmCAJyeXs0kBGYgHs2jKknGkjxSt7nR
Z+js6mnqw19jzzqtdrcsrrgRgtg7oig2qWoYZ02Z5i5773xVOq14Ir1PzTGPIQmw43M0Y4AMNfu2
e8IRWQ0pZeXLYkkLzsohug95fMwdlK0yaBQLujF93oIJBnw/8jJwG5YWFL+WAJyik3d5AQoo49bC
YnRo3rB21r25MiKeTCosJQoL8GWWqtb53YsJNaWeJlhfjkaFSYf/6SgN7FNDKMnq1XIwlo2QaAtg
s6jWPiUw8OnNUcD9q5Ovfifbb2KWohk6EyiuTCUk1isGtqXuEisAr7tgEHFAqC6bwv2z35czF0s7
QPC4Y2ScBmQgLBm7HyIknrNkdm2VaNG0KvXoRe1gtBh2vLt2pJdLRPQJZSw71sWbXz8mY1/1GHHC
Dr3Q3o6VgGi1dbgDnrJ+JKBt67cmdxk6L+Ctw77ssT+qkl7pSjTvGzEnDWfRXmXgLT7EA1k6GJgO
adlnnH4bLcmnH2WYorsMz86iTqaCxIZBEKxZ5Vb738gRd/cHP8qg1YZcVBGT/WSN/nL5darEuOoJ
1n3hhyCZDSJpmlbcprswEcEHB/db6hf7wWUx02zxA0I2MRQcrseKhVemgp+M5UJTSr1RiGD7VyNz
E1PWg73AZJrBbKq+DPh048rEXqRjZFKeh+Kgc3CMlpQDrThqLHlINVfsCux7mLiMieS53vYvYyXJ
LdbQmby3N6tabyoKUp5GODEHrgRqnXv8KG+iziNiLAz11YBAR5SCdyYShxG+h6NoPyuvWDSBo2R5
UMV7V81cDo+MTWtxFscqUqrF5qpqhLEBEyTPrTYvvbI0KJFGr6FNpLfJPOuwxRQMiunrhrhIkvRJ
kyKwEN2HFF7Iwz3IHk+NdfYmAk5B45ZQgT3QfA7c0N7aBK5Twz0gTKwf38ogdXfftuUWJART/k+V
d+z8spmQkEw/JtiBTIdBcV3sj/EsNP+exVuXNr5Q0jiEz8m4E//93of2cJh1ys/L2M+K/kHRPfZN
onY6yGBD76uo1k4g6i/QEGbtpeA3/KHaMzfgPec8aQQkP7kb3lL71rKirKRjTt5IwR+5lIzWiMUL
GvTs50nw2QO8PAJHoR7Iz9knGuSNJDUBFyPP2db69HMg6g8mSNNhgJcMFBLyhcqhAxPpkCR8jzWO
II6UPuOKRI156wVUCaoVvAnNnyvpCYGphaBMsn5NWCl7e5rflnhVCglCNw5zdYloaD8RZeq0juFR
mPJfejYjcknCWphBWNHeDwGto2SF2Dz0fmEyp+kwnp7tnR7hbNNYzdLWCuT+7FYtrUSXBroukCOB
p646L78neyE7pbxswgI1oWLkLwRt1x0C3hbgenjzxhRsYKr7xMF8/da/0ft6ZH5p4f5r/mJDBxJg
8sjtwm5JXICijtbBLM5+iT0EabUwdCGUOhVIWyJ5gOQZlSfSfdIgwThF0OgYFD78ow/WwtJF97NL
Vs++CdVtffi/SKPDmfIc5ZbR1F8k3I/GW95RMSTJR4cGgZzuM1lzyMrR36FWWMaVg2AsJ6toOYlH
OHHMIAv0KawKpxtDqnslhz0A0ohFoXWZn8ciOpQ/vk2s8VbOAL5d6Bf3oe4nfoIgMrRarFFCXgdE
ekGCM2h4uSiRCnP6d3DlEoObQ2O6NjdCnbcFeMXEFNvO++3UvXiR1Fq1+BmyBsn9XGlvRjZL2brr
WCBGoBd28L9XrurpsRnn0Gp2bHqRmBgV3ZtYk0Cpt1AQcS5CUazmw3uJDXtpB99xAHOUFetYWyiC
oRKWaSpiYdGUY1OBlcHXcLpk72zZlw/eW6cB3kq9eRzDRCq4Js2V9FAJYHXLzWlyPD4mrfiXK9cH
zSQpp4yZeCYJ5wCfUwqWL23f5En7s0NvIfIe4zr1AaRaHE/Lf25oVfG9EjZjnP0pDjynkBRU3AIa
bFn0MfGhP09/upl7gvGSrfB7uvmrs2MeXyMtvCVEQk4A+km19xW7d/e+NZ6QpqaUWNCeaUF2LcUt
70+DEyqQPkmKCiR3sTfGomukrlwxpic2SPR2ssntfGrCfhYIqQtS9X/o8XMHMo27XYu+Dke92I2Q
bJsYrfwffQtRrr6xHBhrm0DPW2HQLNQ2i5n/gwFYQ84anwmXHRbXD02j1Y158eWaQ4zlJPfK0B2Y
MEA54gMyaHQD3QQIN7IVbBObCCjKa3wPOS/GjurUe8kA4ZJHYScBrF9FkyZDYTs/lFgIyifEbBpK
HNxYtSHC+hrsZtH2iOoR79MItUH/2dxKSS/wMfX4vx+LLU/0pJthrtiRQ6n+jUAasr5823g1gBJo
GcddtYQaQ+U8s/Qqld3rqy3PAEBQOsF+NMgTPrbLo7zzxDXFvHpjIc5NCHVO1zJ12TIBJu3ye5Xv
862607r5DhjElC0hkwOI4zrCQg/y9GHrLX56cA5wbXEH2fdQtB7IawsOqXkBiIZ1xTJfUQ9UFFA/
u2h5kt14cOEDA37B2y8MWidj8WaG0b8PhUi25mnVEjEO6UOQtea5yEUTHUddo2rC86wgOJCv3P22
PMRpLGe2xhM0LFXhnB+mULS0rgt1Esl3g1EX8zyrXhX2u5DvAwxoWOlq571+jZj9bVbL27zRHPsP
FB72gt1D5oLIwwMvWQAs897E1RP1O74ntZSNEHuOQ/x4jigpHXzhRZDVLvujQ+/9SdhZcrndfg4e
tNZFJ/tmfCWYDLnbX4zE2GZCsXk1E4Lawd8EKgg2FmKEvFk7vk9wdMKbKchVuVWmhDIdDgBFTm3p
LI01GmR0ln6638Jv/7SSD7bZwUjfZiqsqzeOFUSdagjLMEgBNHmxB6j0WL9/Nq/poRQk0v5F9auf
iT9F5rHAuN6FMRwV7uakw+9rgM8hct4x5yzgTT2vkAN0QlI3Oav3oAxkEkZ+vR4tGue5ou8ba/FH
tUzzod8F1CKvjT8wFLqVcYIhKW5L6a7fkU5HCuINJ3u8Gi6IERjkOoVB6tRrP11tSzSYV4IaOPaP
Qanz/yd2Pb5QZujEl/gh3uXLv+7AksEYskLujv/o08wNbJYoIvbOfQEiD3zZA1P09qogEZfDYgwD
00BohVFqRxuj8xvtqOu7yj30BSZhkVacOVh+Y0pZd/F9iHkVU9974nLw32Qe7XmJQ4TGV0qD3f6d
KgbcJnNAkw8THmiYyTkHnMEIEslrXSJhqpJHS9fMWQ2e1DI1zAoHNhtegBSEt/5xpS91V/JCisAP
m/wxBEIasS+MZbATPiBPXvPpRXaUm9ieCULNOUPHEQX+ie+gdTRP++7pZ7QA0F+sMrBCDBC69ie8
RW4da0S8Sm0jXP9W7wEE5Ki29bfvg2uSsNSN3cV0VgIz0eEbHeF1s11iuTEOA3SQit1iF43Ftstn
T4edpPbfY9yhu1ZWNx47lbjqRF6x/JFDuuUbu4hGwLQBeFOOX0qrHM8yqk8l3Y8ONF1n57WV33ne
MDnM2sjDjDx4BJYK9RGiHrzbd3yt8ktk59lACWX5Jp6dz4JuxP+0FS+Rvawvsd1vmXsTAcAjeP1i
NA5MgJP7/ASykTBdlINkKwXbDzvEJIOXuudCLCpvIKmIu6f7bBdfaKzbYX0I+OoULoEnHn6ElpeM
HgUnGEBozSkyowkYbzd3bZGwBgYZ8rLNQHOn2uxeEbn47ET+O5SANfgIm7de+vjwOE15HZo7sCOi
zgCJYKDKqgtaN0nerrRzKRj+idmvP9iN5hh/8PqYMK6ofihmxEdOCtBHqc9X8YMyv548zRIXaTUA
Cc+e1v8ygiKhi/yO0Z79uQSC7xSIDo5Hbp2oQSVrwf2RWW1MMa3HBILL/MKKDX8p3EqDPAjdh50j
xTkRUu3/VcG6DX/lceYB+py4eHg5VVYS+jlfAjyeR/cA2O+I0qkWIO7D/OWEd5L2kWVXm0o2Vk8+
3vtZHxDH+Q8pUEIeMYqFMQM1eF/PSgYYb/o0hrTqyLsJe5deg7jhdV30Jdx6Lhkz+DOfdyrCQFDz
vFpieo6uEYNKWC2goDRp/JadBcwKuqoHwNVjHakkOaUF9sFJfh1gXmDuk9NeWNvjnPW8WCWSgCb3
SjJUeSEg1AsxhmQwGuMFEWa6BuQ+9YG7VXoeexvaYpTzEW71EGBtT4hV2tEuJ5yAjysoR+kKPPSx
eBYdJkukppueKlj/XMUj3who3I5GF79v9ha+Mx9CtLUT1qnXZutR3dfjICWgln6TivGtHq/sjKE3
+a0TtgaC5ptWBZndNTwt3QBSBkWSIil+45FicOFMsIlRQVi4v/ystKf05+oVkuO7g03yoC83VhBf
D37ikLPEQPQNzRxVRu0lEjogubz5Bdx5bBtKeuKBXj6eFnxrN6DNdg14XKYLj8rNRB9Zx6ZCyiW2
6X3+8Lc1oMzTJVDAbRc+09BxQHlQBCrFOUaT4kophp3NseGz+ylEqAgA1KzG8P0FHOFe7+ClIkWQ
fcbWPbJneS1ZILt0SZLcAEyWN50ccGAO2UL0cFdSLXjCmKFyNQX1o/V8vH0orvOodthsv66wzagv
9S9sd+X6FcqaG8lStZFUXSTn9SvfCUmYl88KhEprJ2tN+LPjr+aSU63QP67pZiiIWLFP1jbxOsgY
UJXfRn9PQbdXOMIdG+9G8//SNzvU8XMo4a1LaIFAvM7gHSQD6LUNQ0elYpAtxH9x/T/F5XWPdaNW
GRL9ZUgO3PyuN6bbbXT/3K/2/bnz3HmOZJcOaaFPu8uKBiEGYapKGP7/MPxGDU6p/jyoOWg2xcml
7/GSChniiD4bz4pxwnfgKwVuPRcbkZD4WG3uFROB34lUroTSpmXcYSZ/2Fo9h7sAj1v7FWRln2Wy
DnaWLArWhDj/XTl2H7lFLDlEn9LJSQxx/DaAvr43dmI+4svCNCyV1kT6wpiJLO7aFO4WorHO70+c
ZAdgUHdURA3TCHY29YBmZiv8XjnsLQqyr8HN68Wsh4YIS4qWh58Oxt25dO/yZANMzs+L3WXrSpw6
lAVoBjMvOVj4ISfoGLDpYAf+Ua1Rgkzk/cRhUiAfSreBz/Txa5a7r3+jVbcb9u9U6h8j3M9jE7IJ
hB9Y9SfhMu/4lGUeWjKwkgclbYn4nHO7B+9RqxJOM0q/JgGGZv7gTVLfI6SV+QCaUp+ebTxkJrrk
WdCz6J/agRFp+Sr3N4hwVe7LiUkqoYJpMtXgYzF6FzT0tGsB6d1dM9IxN0sKyv/AG+pNPl/W8icw
vSOXhfez0f66VxKG16cnZlPRXK8JgaMM2FoDqZY9/MMG1PXir/Uf8n3uOh2g5cuAuRnZA1r+8Hvj
Ozsc/W62s7H1LMP5P4qObG/rQD++CZJN6amv2NZsSVvaI/kVUSroPmA7UhnMTzwEHxoUfzYdQO5W
R5Z5ypqJUd1P6XXAM/bEWeTWHm61gR2WKa1aBqq2e4MUQmy1GrKLufsVGiJ4N0gyz/A5BwP8jRFC
q/GXZgwwc+jBjBlQ3TJwtO38PvuCMKJXYis7+QEweMSgtqnCbwqZkCB0Ro46fv7h6ph+2VKaBI6J
vfZuByFlVy9TUXUi9i0oQb8VrxWTi4Xgvtw2Otmnvcoo5MBXkUyLJlKw7UNIBQRcJy/Q+Zl/g9M+
UEh3nC+wykVtVG+PPETKpv/L51BAuKdNKxmanXhpQHmrDH7G1x3GnDac668nFW81EecHgAR1/jS1
vVrCEymMlxUbY0lQmhXn7jt5KA3JzNviU30YhkgSgQK0EnHrrkHI7VWhq/vbH+5D+oG0XBPDJxcv
0AqmB4q8GyY9g1v3HhptFot0zqdfxWmxeK995HUvRxQ7c+oVUU7bxXw57OqR3mW5Jot7RnMKDT/5
pXTZSaXEMt+tABE4t61pYaXtTTFbfI3n2Z6EegF6yacgSe01hgMOaNaYKTO3ojRP/idokwLgqJ/g
jc2KmgaRRI8CLaO30GzJI2AuEeKON1Va0SV9HRKhUutaLDNx4+b+Uy64JF30sxKlvcS70JTHF2A2
CFXAWhYP+8HpRs8JMtxBH0QhokkPv8ffJ2KsD/atulPhAG9iFzhg9w9tIDCdIdzUH0zchily53k0
LPJoCo/OAJTmB8qtS9evygtdLk0eVEfuWUIQMgG9ay/sOZYSc7SQcNb/2gY1FSNWqo11Ad+VJX/v
R+aMOexUqQ/FHq9zhv/QRZ/EJKBoxuD5SYD6ndKBvqYPyvThpzfblnNa8GklSw7+d6wd8nGvjtpD
nOOkohNgpls9zzfeNJUuDgFeZJJRzTg+7f0Ltt6+kumjMWrhyHlGidKAbeDI05tCEussO+seeJaE
+2kCGtUErZq+9JteFHMmGQocZH0rXisC7A6UshOcDQgWzyLVv7nC0uxDZN7tjdswUiG4iawQNbkw
+rTCKfQI+2efsQxG5ewq1kt/Q+hrhSYGFKNRCxvGr/UpLldZHvr7dbh/WzOGeH/VK0JFdhk8St0e
pQ5bwH2XHLRIaFx2EwRS4ncO9HIlxGTr4f1qsw7GLPxsARVZN/8kknVzB4r/Ap6ELC5U6Hj6xPdw
vtqAQ89vZ0PyYDDcytEwotd6me/jjskyMuMRcJN274ylgK8YM2b/LwOaIRpQqiFZk/FzRzNift0P
ak00HvBZWASe6dta/fL5RLkBz+sLCJ61aElmfm14IaYoUnmdSp0bu5+zLTpDEqjMWWoe6XBLH17g
1E9zfPX89eDvTiJ/FGy5LIWWOpkomvp+qs+6F8zc7N/38s0y1JVi+J2bsThonWRjxCKdY+apCs90
DTPx++hUbYlx+B9GFZPBMKvHQxAq+56KWei9XBswwQYQZE6b9XeCyx8PHoU3nrMbMa2/yC8RjRTE
GvIV10fYqCU9vjSzBMAkFQ1OflnvyY3JXsGyNIUePGrzSq9q/cxLL5E/2UEy9+oY/SxITK4reQxw
AcZQ2j8Y3LaNF11L55Pf4KrEjau9vJTfoUYWUymouWp/HECP+7+153JWfuwoVsnse5tBCP8QQB0T
DWw9tPIQuut4xGzOfvXneeLdUCWpwtojvVAPzCas6N1MNVYm4vzqHzxpTDgH87FFtqHR1R9TBsgy
VaWzMeRcc3cIMsX4Wsao7IAyDjtQAV0E0qwbYrO7bP+/XfXB6Twc9H5cuq3NEkTnylxyMtx/Ieam
Gk8BgE/pUtTSMvLukcMcMUiOW54l5JNZ7YXQL7mODP3o24Sk44yCCGBN63VrQhxPmRI1Hx5cdGjF
KLNKVtZ/Zlp4UFSMDLeCFtNEbHNpagu2+RjoYTust4pVvPa75DfcS3dKfMQGlgaf16gfCoCpplCV
eQ8cdB+4pXJ/OeutUCRF6Ez/A4X+0KR4r95FYKk2GoN9nF20Kf5qEQXkWfReLxPAykDTI60i2/kc
AksK7CtxswHS3lfOEtogAvd4NugJrsen1F0JX9uKoPgHPLfj7NT1GcqwGgG08dKoRLBuXyAoMXU/
TJNIwBHGcrr1O0GU0nL0Z9ZkPueySs6B/FdtchTR7W5a+gwSc+31mDReSjzPw69a9Gl3jcYwC1tB
GAQ7fE/s2g0pciV8VMTFQxG+vbtvegAW2gdF2anMp9LjUe4wMSW4aT6zukeFn8AT2yKtAf1RIH9Z
40+cYlbVJ/JB8feiN/paBhxAmUiStmUirixV1/cYUkJ+tw8Ud5dJDRvR5ZRuUWWidZU3/OoZnje1
xr4At/La/jxsAV0oX8PWGXyGmXOHDhTqZYCzzfEYiyL5G2EvdLHcR4CUhHrRevnTR8iiI7lVKBYD
RTN7KLCyYCK3Ogae3JFY7uyhqFwIfAk3P0CHwNgD2pdkJw4b3R9EMT3SrLYzU+yZ1s65SQA+uzX/
eTJfIz1Q0h6v2D9O4xlnU1gEkoBvwnxSbMGyJpywh8B8RlfA3O5TNh2MnrOg5No6oW0RMAu+2QPn
I93+hb9bbPmb2TtVnexoT4th/US1hhM3X+2Wij8Jv+gOXpnebuhhUdSwoSfoUSgv3xFgaVdXQjOr
CMqFdSMls1qCcPqCqTJyjv7QOY53ofBwxFd467a5mbKjUQ2OykkgsMTWiIRRmtp2AyGGnc1HJZEd
am0WKVxT2z/iR0x2XrC/V/Fb3hSg2SBYUYHFP5KNDy0+PKbgjO6jq3vjMr79QjpSkI0vcKzChKWb
F1nyKvpjefvtil+DCQxa2eBacJYe15qXFKS+8pO73mwBJ+5/fQE/ckK9JeDytDomHCdlJiy8QceV
X9AfFpp3M1/08lVdg/plCNYB0Mrei1Hs911/3VaWyun6lTsyDmnZOr79vv7OvJDQT7OKBoK3Dd55
VtUUliSDL58nmnP+UFOPsK2nTfbQRY5Qkwbp8CZibYqWExLOXAvLouHHF/EK9B2a3pGcujQotJBt
mu8qDKyi5KJx51SHi5IDjnVer4xKuVTPy2ZMdLXmK3nej+iCVByFuWwF7XQA5ZXXQsic3v5rlgJ5
XsbFrPmC7qsD1J5I5d9Hhw8yyXxUYnj3QG/X1MfuGc0XBNfYRTJm5tTmrWvzlNoQZRheFiT4w2ep
kfgjkDW4sFjYUJIpQmK97jirNZfh9BZM+zs4rAPpH3T5Nz6/iTA1hr48hRBhnf9AXACpCq4HIFFD
EI/VMoHYsrB2usZ53u5wCeVaaYqfVzo4EiZD6lQ/KssB78sVzBcnQXPi7dfdIWi3OP9/4uqNcgpr
d34A0gaakZcRIKkKRsRzuvH13xItJM9OMFUaDVQsLJdJBynLEg/KHwQIA9UkWKup1vlUE/Bw4vxn
LQkQ24oByngkV5GdI3G+19t6SqpWWAHZLiceoqIyEpELcY0Nv76O+qGSdFXUqtNODHvAv8D4446G
0N11vZgdA/cBYg/KJI2E31vqbfsfOfhXBfUxc3Hos2cwdjO8+5a/SKgU6rjxnmjfHg/1GwxouIE2
k48oinDY6XiF8Wm/UHmZoY2P76gPdYHeEdEYYlCex3VVkW4Zn/4dw+1qLBq6ugyzFgixt7AqlWSV
xn3B8wQ/Ht+ixY2O0wNVfbuAGGIBbA8wFVFwfj1HsLVKjO+AaaQX0ic6uil8zQAQ35Lq8vefKPXn
lKX9LnJmqY5p4XxyAa8lYPQjFZImpdGdYw74C3wVBUEDcb6Wd5hV3mom7PysXe3jmKFaA0oVre+/
RAcPNKBel7wvvI6uqK24t2kwtDaztJErcGChg4XA37KNnVV/PcGQXjCpoEpLV0eejZhuBs8T6uns
Bei4Rfdn6cbO65wpNmOcavfRcYKcax/3CvJHjWi1eKcUcB1UziC+eZ2iCnCiUAgSt+Aj+rvVQCxF
OabKJGMet8hllro9iPkqNL7+pCNSHvOQrny5h9ZNYqV2L3eHk66SUvetSGTJN1uNh5qAKPHLewoK
HsXUyf38kb02vWWTmML+lkUT8JY+S077opj6ckL3NxdiU+8reW0FqFQA2CFDJC4mGKNIf9dtwzik
GAqKHDHZSssWd+kODAuMt84jtIJWtCpEAQ4oGkHpBuUh7ekKR+pBi+SZnN7/dVyXxKlReBW6oFed
hOWO+7BuHtGgAP1KUHx0+sIYHYO/nmLY7F5VP0/eAhmKRlf+hUvaqy2dgC0+/j+UTYhdJvsMH2CF
UW/p3e+6FTM0WF3ugrNGTB+UJxHtXejYqrsT4RCdM0aaj67UXITek+Hp+Fd+gPfeqXU0yKImCiYK
455KhKD+jWcwIa1Y2aR8lKmJ/NSntK8TnccouxcOGk1S0wvt/Pyc+vYAtrVdPT3HKYpTgrM/RWHn
371I0VAI/aSHnmGSiY2XxZpl4/kQsEU3XlrhdnqnQDwrujuHu930j8li1R4Hx3ssN8ykZuLAO7ug
jDjBPmq2mvnT1a962ufHS8ljPURVMODLNKgdK6S4qMxgXnJB1lGsI0iHOsc2puYD1JBzukLs/yR3
J2z3wZCE1WUv6iNy1+9mp1otrM33Pgpj1vv9c47+w3VqvSJ6z/m5CEQ+nxLJJwh0PzVKDyf/QWa7
8w531P27zRnyAIbrv0H7R2dQG/aM+QsehU3SxQAOyyyg5putHcefSUK4a49ikr7f1QeSRkiLvDnz
tLWf6cCu5Zp1+ewP6AS1OO/3xhUUs/rxv/VVvbwS0Wsmq4o73koATGyVwSq97aKoSVo0cxhZExce
XEm5/ASK4S0TuoV9pOBT3D3pUvn+jhGEgSARSDx5S1QXqVAp6iVgMgMvJ6JBfdaAu9aw9hOxO7Vh
qDtMcMTB9U1v+5uiWVkz7qeHMunsZ7yT6TenVRoAeP/ZCFVJrb+LJ6qr893gzZj9fUD2+SAqI/Dz
/1rT8n0G6CEEFJDApsSAeZi8Z2qayKbj9EYX62uwfhPUvEeCr5hIwh3spLQMejicLRuUo2xpGvVo
kwfzb0GnyqZW+xmPIRnPSqGHnWZHi0ORrLgZ7ydEQ+Dfz1LYLy8BnM7zVmHJA3zpLNSuwhRIi4iY
UW9DiH1VNZp06VXkpL8akaFy0OOaZzEuyqlaKs0t/N+aigbjPvYzW9owA97EebDM/jM48U/p2Nor
XxDp8PHDzfFs2i9PH8J/GQeTaqPmhWJV4dcT7ByivGIDsxf1dVr5P/tFU9FWbHOmvVXTnfXq/dIs
pyLcW5okrs88ZH0+uXqXKUJpsJ7K6yy1OtfLUpGSR9pPWUlY+05Uc0Y51mNizYePIUTqTxGUq5NK
7sRt30Hmm6v3sHGSaJ0HAxAlKDD7Tliw+1NnYBOTJ1jR3giqVPIJDoG+nIpKcLQtp4weypDx2KFz
gKCahiAIxEARKzoDGdEwf7kq8+BCZ/TbA5f/GRRHTdYG/cS6T/MiT2ZqovTpdJkphFzOsI9Fzh2S
sqRO3yXsds9DXbtkED27QgRg+NiyCurUyfK/v6y4+QdOZhM9n+WaXASBUgod8CJ/Rm+Ntnj1f7cw
oobVKzJkqQ1/L9x9np40YeMZX0T/LI9Te9Cyhx+cw8anQQyKMKade1YUCj2iI6mCqaDOkgsa2tZY
Hu1FSI26hoAy8hCEpo3Er8WUKlaSZ+BAtiWL66brLMCK/OJuT1tbMGjjnXWuZqQ/eo2mcyWxKpSA
v0t3XOGX2MmzdDYx4pkLTy4rYk9hDDHGU0A/8MtghzVe4fFRmco7RdTkZYLBNoDsXHzCXUO3rXR9
XgxPhSp5g2bAIXmjkNyrxbT4aCSqz0VIqFBiv+rtqmo9MsTfxYSPtChzxY+wLsol/HKWGo6tgqvY
WynoQBJH8pDq5Yo6zGM7++walgtBko1P9LRpJqJZv54Zf3rx7at7SVpfuBAWuiG87nC1AYBNH04t
LDzLUMB4SBtuvtSItrXtxS1TpLAAExTYqoL1KB2RS25MC69NVYEc6ds807ADfhxXlndOOlIAlatg
OSPz1Ah8hKU0L1ss1LzDf5cz3hcjV05LA1WZBd3Y6R80I7rG4zDN+WnwtZDLZNww5GC5uzaIa6Va
0lc3fL0s9tltjgxadHKPMlEwyIH+Cj7STrzHI7cL2y1UpImmAEh+X5mJ55Kk+1E8v5NDbptDQ+JC
9yKpheTsyjmweVW+Qf5+U11RFNZ87uDHC7/OLGl3zxf7xkH0Q1gPn7tLgvIvW9n4DEhM08pV5vxm
XdxLdJ9vro57SSE6/7e1kM3Gq81nxBCahb69SsKEvsXAUvoEJ6TJ4Bmrfu2kV+aodimiTKd+5gKn
Zcd1fHFhqbNiJPLTsoxkJATwZGIJhIQtw7VDNGM14Yjh0qobNFf/P4BG0KEz1crNEbwBZZq2OEEo
lmOwZUk39u+VNdvn/iL86hdJzq/CapXPQTTxCRAwYWVfJ+XkMciqntHbFDvKqHSly+uQ2TUmOSLv
P4bAwHahAqR3fEMkzJn5ZkJtBfWaALMSC21UzfU17GZn94WaDvezfCgibBRa0gJVunCbu3lGcqv6
2hJWEXOvwYwFTsznuzxsY9f8glK17gVS8ZYOfguqbWe0zPmgM+lH0JoWHAqohwX8MKxuv/v/rR9R
a5ilVUuW/cLOHMkV4IriAUPXJKQ8f+J22jtto8vr4q65UKbc23rN8zwyn1m3sBEBWKB28xUIIrA6
wRnDaXVtKzymilW4XO7gZ6pSbvV/MYVS3C2cXiluio0jgB+Q019A5lzV+y+bWBBg//L3BAjgPMzh
9N4e+n2GGoN1IsHzBzVNRWgZln60fmwEG1wjgah2Hbapxy5mP0Kl6Uv+tcFQOA0ajW9l445sn+Cy
xVmWydZocJeSXeyhD/bMcpw6l8Q5lhJXxfZ1J0JQkaAFMrqhME5nCf2ML+DvW22kIhDvQcNZfzUW
Dv2+LZsyn87uENrbcdtnfFbJb8lVmc+4Iq47mZd0pwWEIHVZMmkdiKgAuvaR4kqJS506zhff+KrS
hiHaPAv9S+gfh2jv0/2f+EF4c/GAwsqeQLGTyJMvOqPDiNlMd4JXwgmD8r2G0LCzfRsreq62jkGB
MHF3yRQstQutrkef1fhACshvvCtxO5rSN7CX5+vax8sWvpwUFdspWr/qc1OTZXDQmS/ltajX5f5r
aV3gSKD9PVQQ0yhh4ZJXadBGA6kqGCAolmR7waJtd7d0uV01I6F8qqZ7vrzvNkuSN5dOiZGG392o
V77cZhie/cCsE8+KYgA1HmmkFrNHGtYZOxZcdAQMNnraDzg7Dyt+j46DRc5B0TjLF27Fk8AofRhp
1EEDV2RwsnIqsqTlC7Qn2kmDNbcv6/RFlAGbHQGunfY6JbG2OlGVzKOqPadDs9khsWJYW0/m167n
nfax+etugqaXPa/VT4rFq+igLzmL1/XQx1q99IZvegTnFyE2KqjCYXfxKzkM6p0y5SGFFADvWJrd
BzLfrOIBfql+rX7W70p/1yP35CrGdVyhg5PqbB0QsOwkEacBdZdKufUiQPEvAVlB0WDi8QgnRdyb
BqPq/FAbxDJ2g/7s1rVPZdZ0LN4CklL7WPBbzAbvki913VDPeriJX9G4UWDszstkSk/D5ck30M5M
EaAHb+/t6YLdz+RdPPwAWTfUuDoZGm4Vr822DfhKNGBE2gvGZ5Y56ASzNkDLo0I0nXQZLX9JXm9K
e4oUqhlrGEyCsMsoAC4tGhCv4q/5MpVpLvJvQ41toXkuslDk9fEcwKeO6FvhYjz5lpzklMqm4pDW
8dVfb8q7GoFlYKJ6z7QPIqj92el7XRL+YQZnVW1xRE+fJs8/WhedIY/PIyzqWqPFnovw6Z12H3uj
NH1l7SgdtDokuh7gegkPwLVlFXGnGhlnkafT0irNv6ckzCc3rNFVRxBXoS9OsDo8EbjkQyvnK5++
JH9233JSB70Gqp66lSLp99F2UwsMElYK4sqdEQkWAW2tnYWwqpVekMlQTaYvfMmFOPy324rSEu0n
YJsDXsLoVtIEgAYlP1ThbN4uyd3zcI2YUqZez0ncDcWCAuSY/JIwypfnUsjOJmC+R+kZQxfV7NtB
P8ptN+3L9lNd/VzZ9vNFDhNzpXHQVRgGtJPlXAwoiVHwkseaj/AWE5Qn6m+YUVWnAnJlgM3X4kwA
R5Cwamwu/F1pmVW3np7p/jGe9ly2dpyhJyEMqqUscR9JpbX7lK4SgIhmNKWF4/jyGEKQhnGvt4ni
mx9A5Tgb65GShEHKF1bOP8/WYe1Ih79QS5oUYoDNxKtkFzkW6DexR+x02esben/5S/Lfbf5N1ZxY
74qO95sjKItMkuag1kzEsQCnfHIVH/LHSyv8HEZhrjW7OTDJKvzw6Lb4KeFGdoupNLxQPsvBwEk+
30l0VtbhgAqWcqJCZ70grxWbXA8OwE9e7/IUfNuU7ZvB0Sk4r6pEwikj2GdEl0d6Gv3jb7VfPfdx
VN0hFXtEDsUJeWJzorRQ1S4WWgp44A+pmWFd4vZ0jY672utmUL+9btJlRJU/hip5KKQ6HOqREBpY
SM/zsaLoomnpgkV3rDKGdEM+mEF1LE0X41esdxwBaZdQHG/kMoa4PpZXGsgxFM+DQf8TORjzmiNP
uVdycdUutGps4zwswpNmVQkG5dat/Q2iG9zmLvDsAgb1o58BeCu9kGeYptnOaxyk+9fs6MHugVEi
MMzHedDFO36bJXOsz91fUPYEicVCpFlnSqefd/rZH3mJ9ANO1lC+hu2UNxVtzTOUCNvIMQFF6dZ5
wzvEuXGeW58vtEHI6X/iYiAM1pj4RSJ4AprUaVFoFN9oc0W22inPWKmGAtz9YYVvnnH+1tb8QIzb
0Qmma9mXc6jfRkNiPrG6didZvqU3v2Z2O6ig8SFbHCjSC3GDeBGUVDlI9dpGGnMfHxhCpEAsXp15
8jluGyiCACYSWgmFI75cSDKBmp/pmH9OSkynoq4hNWwUpoYNRQ6GuOTbpqwt0YtEoGqnwkUJco51
ran6Sqc/KHixDxtDTVidiwfJj/bg6TW4hO/BKJnR13JurPs41rrJ6RaNdq9pHHteUaX3qFLkGM4p
gJkYZR/wInqBzVBPzX1OeWEuGuZF0XHt5xQT3z1ZnuFiTJbjxefkRZhHQn2IQ2r/fTsEnFB4JCM7
C0I3oDcjQwfrsVcxUulPJGQ+XeQRMlaBpOxMyX64zi7ehK3ZPNv6U7KWU0nzfQE3mcXkL/pBmdX3
Kctw5QSdXBxOy7zDeITWJ0pXfyP/sgvYNHAzsasfWrEPIJIP494Q8/CsWV7Tu8DBzrLIkMUDvwSu
TbXxh+hFu5CBvSXIyoua+dgR2hAJpnR4Dv2TIh1SEBPeDZas9BR27IX2ry1fFM/Cw8zH27dKt8Zc
FCxn9gGFmUEkOJ7nSPFlRG6WsghwEQSvbYE3c6dAc6mU59I9TEtSuMD8CYazSIqVEWTzTmFOb7Vq
IhkvL5ErLQTDnO3B6TSJlqIlw2GmQezHEoMt0gu/853cxTRxPbp4LQTRa+o7Q9X5T7xryxZT3FJw
olYGWY/jyAeNxOYrLxngYGed3GpENJCzA/ZGMUMCMZ09IECy6LDiJG9fWzBgKIf3NHP50BvS3lCW
5ZGMLu5gbHafHtQBNCXgZ89ZNoiwQKcE3cizhY/7bM0fNsaYjrF+h5BRNSwR3a36DbFu6ZSa7D0/
YlUNuSANbcg0K+xqFY93M8O4W+MHyr/nlvGf7gsNmQBqcm/wQJeRJvzK1Uc6gHjlwpBFdK1OuduC
oZYPP9oDF5HKrl1MP1HvJNBlkcxzZCvqrTWX0tgFmvjwTGD/m92Iep4ye3xZFmV+/acMcBX7Z9AQ
yVggdX3TQiuPzqsSDkNKG4Ce+QAPuF3tUAkg35ox8kd6UP188L6ZlPl48dk39j8PzpmZK8T17Clj
Lw2hlJU3vKMhZcExjJ9dfeFXIN6uKGD26tsgW9m2gzic7x+2zDmvt1muu+VnVMal9q2lgwFXo4h2
eUg9VtpY2VXWFb1S8DCdzyjUT6+NY05k7QQ0NP/+LbICUSQlyP5FiszmgicVAVWRMCiOfY6tT/f2
knupy1EADB+Xeho/Gc31aKERsDnXo4p0UF665F0tfWUTBhdUSMb7FaL6EGUNdL4YKkrH2ludNc4E
zlWsvccspeh1oqpW8gq43ieFY3mKHNSuAT9Cq/jNvdUhN6G6LSCKeriO3hvMq9uByfnDONjFo5Xc
HuzSboWmXt5DDzrrCkNQC9IsQT6omGiQUahyUFK+HMplN3F0ivrLFI2QnKaBcTwC2NTrdLcZ+bZ5
De+dRrpuXkgosPCRVI4+FYEfrGOGnQRbMHiF60/cLUhHQ94XIBPLmWsHh2X9E0l8XJ901ZbXTSxH
V+8i8DWL2jpUocY0AW8kUO2d6aAwt2f0RSKXgQkfVdLjiSA3traKVZIid2MCGfw8UtdaUhGfGDjN
PEdvXVAWhyW8pM+iHRWmn089h4bYoXNZRH8RYCL8XIYWIG8EfSaBSEYH5bfTyMRmCijOEAKwVoCX
5w7zBjKKKTEZa8Uw7o7nt8X4qTB7QOgD+aeUVCbc1SjkS1a7RxHaKErCnDOpqEYWVNUO+DSEZx5s
hT6sA3wFRmq1bRH6SwfncQeLykoUxz/f5Z6X9j09H8ihkrKxW8iznml+oLYv+f1wMCkcOWBfvpED
hOa2r9CMVwiDY/grflolXbThj3qy3ZcaMgCO9gS8KXHZBncNHl7o0N35a00Y4yc+TR4BnL0/I/ib
6ETAMmV+ISOJIVuadZNSNpNS1CPvBjHrjesUvuG2mhpE6LB8ut7Yp0qMB6NziXpZViC9V9ngL98G
7bd5t37k71IaMDrampakQ9Us//90PxwGHXEVYxsVqSmUx8zD+k9Po0FpBNnUbk6IsyOasUuLSwXF
PefUmY3lWnQYhSmv1h8K1tq8+/7vOgFAXTNXaLfn+dm33rlx3TKKRlxF6kx7e/tZ4H5ACyjFTiA1
dzbUyQLHN0wyvrCC1lE7rRnUZ58REOwipV/b1WdjDekfnGWbBmm64sqABLO2plExEi4NiikTFi3P
09OgHVKJxfmkowzIvVZZ1dmAFuYn+gVP/NtaUxdIqC6KA7HpatlTdlZbBUT6VdcPI+qRhNNrQsQl
uIPKzVeVqo8VL+sznmTngmdc2VEy6Gm9vdibUxa2kCgEISKdc1nrSG7kGL+iQ3O3by7EB1m6cxbT
aA/ZUVxxsS9qCOOjnrnyw6aU5rGkapvp0b1yzHYJ6DEECc1AgkEI6g0mi/CAZiIcqN5h+x5CWQrD
1FJokaGB2LKDyixATXPu/6De/JOqaHdqqEDHsTZlnSnQNIGK7LtNFLAP7ER0zW3Sdx/dWEqT60hN
MnyTelQpHoD00EREWcjNNuKPWo1mkDYq0FK+hLLFKcunNPFotNEeJRTeO9PwqEpjiX9TIPgc1zQZ
RohlxFM5XbLehLSrjBhFU95ZMzHd6rJim7uEUNe6HKnPryAb0gnaFCZ2cBZk3sza4ii+qJSzHTQ/
WnYEtzRuCmLdEkSgr9j/uYDr7IZv/bw6Rbs7r/Hjamw3qdS/6WSKSxot2cOs+G13o2dq3QJV7t13
qxUKHCO9/IZErky8MeB1V0DPtwxtJRDxBd99mO+pTTA6YRhtIeWKsobVl4I6Txn1RgITsp87/nZr
3YJpvq9jSI8xWFh6VsWibTlSAG2Wws6wic5N21pyN9SdIXVMo/s2dBd8zwMGOc7yDdmcirJQ2nlM
82e22NheuOiUXBNBAowohcGoaIZvcA/WVtlyUI48MrLQyRvRto69dnBICLFfgtcy2NAz+0S+Bglx
M2cBp0C5mWpFhReS7siAGeqkDT8yTwFIj1faHnADTbnzsL5EpCI1w4/vCzQMiWZtEqo3MLyjU7W8
cLcTna43/TxdlRvTcF7ijvhp9AdYnz/5E3spfspSDZh/pOukfFp+X+a0e9elRsX2DRtlZejbgISM
gFf+DH/oZgruaov6J+jtkBneYSlQ0lzYL7Jb39Ut5di0NXM4TS+I+ZJIk2JhYZWC46cJU5kubScr
TGr6F5EJyxXbjqeq2iQXJsIcybeay1N/aaZYsFkAZhBlqXEA23ZHx26qrfI70C45nlr/Pyre3g1w
QXghcIlEZuKWDWa8iYXs0AgRpz6tTjcifmLRhjghO0BFo6eAM+Y04qEWhbiN5+dDjcRjBse16CPp
0MdPJO76LIfAkEHe+fmpUp87NybIDW0Z+l56zTdJnLAuu0vdu+E2Os432PgGeFjliI3hYBuUr5e7
DN/IVpFD8wESNYqKC3jed5pgFKFGG3K7vFTQbnnRDl8RcTAPn5vT0VwcvBYgrjhdwsYzCHBUF1o2
Q3IB5xz9DG4jITYXjJ5w0fhaCz3d2/2jJ9c9pfmgDl6SyvoEzf4dxXCVPiqGjvwnpHbClSBAiwN/
14qoLh+pMMWuoBzanx1jQcTDvNdfdqfr98jaMXQe4AoU6lpfjehwP15VjhcsKTrWExjJAqR0hok5
QFSoO/53mxusn7UpfG5/TR/rw9X4aLkUs1lv7MIEa0d4LWd5XQsE1GSvZXdwCs/Uf2CPwoY3yYRS
jMsoRn1+Qu3snLBv4uDqxwnxbSEOUwwbeeIYKoX9jxZpLermiTJJCvZ/pFGD5NjjOjoKlTxaNg/y
mox78QOP6nlPxm/l3Vl+Ju1113dm8EAEWh1u4sGYwSU32e3Ch/Nv2zDGXoEMrgxIW2k7he4bmSh9
QxRBfSerOSUvZylsb0nPQ3AiEuoP9BeAzIvT/RgfO4ThdGQBOMep5hg2km8btA9kj+M0IPXRnxJX
v7ldseoVkrTpLgMNwlXPr/UNvua3wBGXxU0Inx2oOw3vAPlG/38tVZXEeT1hOieB/NYCC52tq6Z+
tBL6A66ue8JwsZe4kowdw3vhE/Cyv4RhIIi4phq62kRAjLpB0P8LHfqzpy+UKDCD5P/VNy6R/E00
xH5YaCLVBMsQf+L7NbdL4+6RC3N2Qioz/9TCuYiRu55OsQ8o/hSWgXeCz7HZkidc1ZPZ4+5dAb8a
mjXho7oOw/uOPETNVRxcJ6ADGS3zNpE442+/oQ6Rqu/aK5lSnzdRFZGskjouFmx1IBFqimUy6LME
IdfCfJtmCuR5oGbptbdvS/d7UeqvGuWsdxOI1o8Wa3Vb1hSrJ4sMnEtO5l7lbzowQ6DtxBGBi2A6
jdcUcyc6/gPPDyWRF3oz6Eu60JlA7mnCn5FgzDqGyX7M5gl2JCMC62XMHevqUN+HmtfTSDv6K+FM
YFLugFHJE8VSAdfUVErW1zPZBJcdvcSisB+95Wfspnxj4+/z/MivSiHlU6IA1XCWkgEP8P5sutFA
t1FKtmxJ2sIjdJONESj7s2Cf6SFqD+Ka0/PA2MgxwjP8IDqrzyFCXDu9h3aNu+If4tc7BLD0XCqj
3gd/znWEhKiEsR+L57e9G/frs4ipGpU7cOCSED7fXsm8LcDhhGzEaoNHqahQ949EScUeBT1rQKhr
ZjK84a8TLOoknrjgwFkMu46/IX5wXNlqyUE+snpVyOli+6XqlXgrmZsl4M98d1GEC/zm20jNJbnW
Xt5kZgMym77sfdQYgKcPsn3mz3OxN1a+Ilfa1eq5F2LwZmGr+/tezj3k39pwPaljpocSJFybck6l
gbT+QeatK2uBxj0Le7JsGvaw+aK+lnREL/8vven+eTWb/knZzVndIRCxnM2XkJHQOmlqzDoHm/NV
yaN66Zb9y5RHudqab38kmGEjpLqxnd2bvirSL3REVDMpRulHoTwIVrPRMGt1RRInxEf5lq4biSAZ
Se4dYV1PX1Iz6a0vL5h+CVFs4U5eC37qwCigy6sRLukDdIGgDLrXe0Wx8UGQ2HDafMag2L5FjRQE
k84FNJgib1boWU9Rif9/ENRMnCbHfU7h6pXIahNq1gwJRoaqsdhF0A4S4o0/2yrtmiRUdYB1pgUr
GUziaYerh1BPz+59S2nvXodX7/iaMexuYtBzLPb8yv0k+3nFjXXkAj7Y3SPLC+Sx4pfg0rK8A6Lb
Qw0XOhzB6NX5GPiYqGM9/qHXvCYTUi86DXuJG/yNfpQzKiNt84wvDK2QBwyUZAmnBtTV8rGinqTY
dh9BIO/gSdRB2Z1lqn9+6T1teswFXB6GtSBpr48toqKlxJwnqgSLAdmiO/YNkglVWrmgPKyiO8uI
URpvdjEpln/DfbP1EHrwtqD+310zb6eLMaSJxkK1TYU/2f54M4JyslI8nlxQVoVJ6MqDRKdJjgGs
5BB59Erl4+LxWBn9QVxs9aVYAB4AIPjHq9h5ctUrsYkkhid1BhRAwQZ7zFH6bp/J5hJfLVhTXphU
vxqC6ms5yQ2T0PC4ctSmGF15R4CYbU5lpWrx+8RzkvtI6LYd4hsZnybOhbdGm3b0enuqFfYmR6EG
g/W0CdzyZ9lsTzYeqR9hBeCXv+/zOaxf++gSVvZFPuOchfGwK4aEm3/WzbGA5BU7Kx67wpUOnsIt
R16UqgOtmz4CFgnc2CFmeYMjy9gXkNBOo3ALN3s3FRUAPP163Sk5Fpm8iv7cgLKhyzlex4KcPshC
/T0Rg3GqHI7wUFKggNmn6bSnr3UmJSq4lPZcLi92sUKEIlnV+rPTJ1WKFAqrk1Cqkq/NjIJK6hMk
2MbTVEWPTsD6+AdhEEjAyoxYYKrMP2xX9Sa+/8jdr7lZFJCfjyxGaSutMwm8NQAMX6YN3a/3irom
aVH7KbMjf5CxX9DsZG/sLS5UrXzQ1fzFofE/hX4vhgV0warClLFaLJ0MaefxuanjiLtbfsdxQQQA
dfdz2bXmxnnMBFGhvMXvBOHjQFyepw/MbcJS/pCmB3swOzNN6pRpNlQrZihEK/0FCVwc1fjvCd4C
NMOwLx8W9zcsZJRO8ET2YFaYvmlSpZRIEwSnH5ofTAwypZErLirgjAHmLQuKLdZHyYRsA/LphGL9
XaTs/E+HH8N/vGuqXd8dgZrMstNtkguXP1f+1E9Vz8pqYxEFmbFjh2GB7ExIN8t4dYqam8rgskuj
CYiLvOl/+0YbGGfeXm/Of2qB3awaqBlivE/nLK2TSL1PKs0NxC6yQBN/Na/tgfJp/hyoRi68jld8
MRn/sSr8YVkzQLLii5WUHh+pVILENNma+gXM00tmJrDeiJNIC6p2vW/Joy17XO5HhyGaXP3WGAHb
dqoUwKC/jsmybmeYAJClESkXoauxsnMHKGdXoNMu0hUnzXcTPpXjbnk4FxV+7c2vpsn0qVBTdbY/
541X0XlsmNRmT/r+3g7nZFmcfT5ahoGY8e2RCGzO1ng5F6bhnWnwnXJYEBwy/vRlDvlKJ3NO8r2A
Od7M7AQFlfKcpMvoRGv7DepYKEkunqCBdwnyNhf3KfFcJAQcYPGLo0bjvUgUpdfFAzPaGCxob5Dv
rUx8LNZzixB0bwaWe7xJBRzSXFM95b9NkVWncMgeUe25Y/CEs5zD2EZ9uOQsntvB1Qb/ygPihOZa
k27tCvVxbGxEQgM6SkUSWe289D7RMtx+uq4DTxz9RHfGgq56AeG5eVhyY4AIDCHElINYWJq7PPUM
i8+kHpt8sZ7rxd3Dx4n7rQlRGpVC9dN8lAt902Cs126fqQzPtxjpD3r88YGufdcUZ0ZTo+/IAN2S
owceqtq62kwOg5P2orStAbldxA9M18VGXSJkKY73bFrTN0lvVE/FQEoVryEehSiPWHtc6A8ui7tT
l/8kL6vOE3hsQfvaUTBJjTtwWMS9qmAwbi0Hfs+2aGeBrNVS1R73UvWMs2zAfdP6qqsEPE7b8rIq
ic6slbkPU4e5B2ggpkeZscG5gDFcvbb1NOIZYLKCfMKdyILHi2UahhFVsQXI2wXzuulo8mT1GoTT
C4cSFHWlSUETaFpGitoOAVGdypmTjSCfe3trgbQZ43426hhWGnId1YPHfTlE7IAtawVpjxQzr5LG
UYkGD8WusbjR4W610w5Q1pg/9o1Ue+ACMXMzU85oxsGPCOkK4Uvnx54UDjGN+2dNADFXZbFglksn
DGaqzouRKEAQt4Q89+Ebjbmgs0W6mPNBw+iQAjR+qZ8r20xOlO6paW8MXIEfnk9OntsnX5Y7pXgQ
N9emifVP3niMm9gxzmv/FtmablCbVBxDnylIStQ265Y5O08f8d90vIrMQJxU2+tvd5ptDmjOYtCb
+buCXarIqYlvm4jPn1oZg41Uaia5PdukBJpanXxdlabdOXf5eo+hVNWF7LcoBxppnn2YQjHBdUbv
+u+CqCDXrxdlcfVo3qSZe+YzWBKLNJFKFuKEgBY0SJkUaQYERrqHKou/OED/eEMMvxMX+bwnPK5L
dXC5WrEGhOvcfuU1FTLrcvKKIAZGZVv8CGLDjM1A2DAeZ3GdXP4M0DnjQKfomgnR/qWgEmWf3UYg
krQlGTnUxgsyLOH3rn6t027klBF8hAbNCh4cryoTxHY2YSgW+6N1/elZTTzXjxTC/1ljXxMlvVXV
AMpv2EeDn7P3vHhqfEJ+MsrR2Xs5BQK2Ljx/4ipNaOFdoNtu1P5aHcCYL8dqaeHAQ8X1QtLDHWKY
TgxY+Z4uNZrSRmLFlGrLxpCnzwVFOKbuP3PnVsNLesJmrN4wOFCF8xz5BbfcJYKG6c53n+ExdGwv
OuqUFKkvadEbHgxxlu9WyCHhkiv9D83b502zPCd95818tXTstLvcv3hqGv8lXFydVnir0djZ2WrT
0u+0/CAh3Ge47Da8bEbsmqJJquFCvU14q2Z7Petg9lwgPRUeICKHP9DLGfYv8iu9O0NTcJnHXMDh
Izy4gyUlDXyhuNUCwb+Tp0nGNFNUDILbX77JdsvKiDsScHSLl/HIiPPVbbdT84eVuYa091DRYX6H
1Ze8ekHqtZVVa/BEeM4lU2uer2wYgDpwbXsIzHbyGjXT5inSAd44LX/wXbN/0qBK04JITw59T9cD
tX4JN26hDLphZhR3JDD+jHLkVJOdWzx+cBmmYDrmXOkHvAPYoNF0LJBE4L6PqJE6Q80yVaoeDfz9
H1hTrFoALEZnB2JZxsQ42vKv8sQsEY6PR1GaKF/Tm1ddnsjVEP1a0IuGqf8RJmKP/7z/jerPezgK
ZvNejdov5221sfLJ//1jW+IBS2cEmcg5eTRpnqzxJaG+bVLvwxHwcYETLFRZLZH2/RCuRPztbx86
mBl8vUvyCmIajnlzEyizL5F/rIQgWYjopJP0E7qOVQlyY109o9wfyo09FjKrbF50X0fQy3nZD3+B
ZExYxFPc26Cnn3eDvtC14MG2T1F4OKcpm8yC0KNA1XeTtQRiHuNFDFEqQmWxf49hCybCwSL22eOL
LRygKXrzlHZDvHUalOJS4lTdnnSGl1dEyRZPwT/37N1Gv/DrdmkFvXrHOSQ3YfiZJG6u0+IGo2tt
BOuuv3eMnRPfw2gSbUOCrzDlBv/SJbfk9KaEk/Ls6nH40FMABxTMcQzZWUNKL1CX/6le9i3uqH4g
bS3RWtAphoJPYtj2BvkOdLYSc8imPB8yyQD8UPkEL2mmApYMlLStp+nXiEk7pfE8BP/ZiLo/OhIs
TIDVe1UNFEWSu3yFoZTolTmNaEmQnzQHrBrPgM0XIJUqbW5ZzjgUXyD6eiPHTek7CXKAa8jVfrgL
8VUL8zVk/H8VAr7AMxa2nCScry4E95gtoxVYvx+9cFwk+I7CRxPg+iHSoWRlixIsYdSjzk1XD8hz
gnHjTnbCs+WSK2wharD0aM7HmOJE8nb7lLZKeMm6xLn8mdONAXxkQQPO/LgLXrlfoYMs/v9y+uas
X6y5I7LrQLJdf+SiIdg866DzSxMaTMovCL7qjX+s3BMnyVgkgr0iv1DGd6uX3hjxuN33GrdPEJut
pkNvmu5pT4j7yxtxvmieA8eWjCfYJzG12aI9DJMOIehfw9ZZhACy2d1SFVCpKu2Dw6BBMnVoEUT/
RCCYKBxeTxz2sUCNARXgYhFtb8sRqgWZ0G8G/7rEVR3Em6uA92EbkwVepmYKswzl/o64CYBu2iOx
D4mQygFZwBkYT5Em1jrl/3X3ApB84mHkHO9pk8sHBL1mp3Zx9NdXVSzHY+CM+kzCxJFUiLoCktwH
tA3JZGCjm8hbuK8lQjRhH5LG4iCminOxHXEAS/cMq6wVGPE2z9RpKHYx6R3UM6/0Dvkj4u89jENh
+a29XYZRK/yIxTdgyscevCiDXCi+qdkOS3ESiByPrv3zQ5uEBHkEUg/zyN9Cf+0rYxbJYZCGjCTA
b9x63qNO1p/Gmjno01vrdpxUq7hn0DERsZ/nye37pE3w/ypd9hf1n/w4urDy2jluagEO3A75ZtEi
aiJ1WKiFrBCyOgxn1yp3TfiVK9EwXwX9Vtxu9mAY1yUq7WNScjHdzBITKb+ERN7ru5+9PY0QWsa4
p/235snZMaJ+jB0ZAGN/V0XaQ3XQBzQH7Au+c6RDd2CtzrO/vIuRe6ziH06gzOr2mmFnZZAlpnvu
qrS4XMo++dwhQJc00riy24BnL+vrYKInGYkTyYlBKFleWT3EcQlBPyf1pw/63bsFbXJjLgyWhRMy
mWxPy/dCAvqG7Mys5+wJMJ8p0o9+C4vC7pyyDw7JIWgwIBGe+T0uS37zVNz+ug6CuEovS6G1F81F
FqJSnxeDmNramy/Eg5a4rkdNzNgLqEgcUOvInRbuViPILO4udmtqsb2ZjETORNcxGgm6qpDOzfDV
K/idz7kw0LeuI8KFdaqwA+hKvZxz0TxAAdJboN1bo0lJvm7z4peEKCSwNy2ls25/KmZT4Wp9eH+m
LQ2yuEBmh34tP6kMupaZS5J0mlVMwt4DWaYwIBHYkmPK/b1k0gpBGi2wVr4J2NugiqYEf9oqcweD
+ztC1v5U1unD77PQv6R1inkJh3PqgcMqRw25TGreCgvEUHdXRDBEl9H4Ext7YRRQRhPRtyRtpSxA
euS5142F4q4Fii28VAP5S1lQUmqPmXuBoGMYDJTLfLjEA9K2Ple6APPr9mTrNxHCIJ/Ft0yPOcsG
cYPJt8Fdbohjlo6hnfKnQYZD29nMeDhZei3EwDWDWsgtOPlj5kt0N98MEQltKgeFwOFD53NfllKZ
0QAewYZvNOAHw8aDToZkwE/cFFqgF1QR6kIbHuQEJ9tgU+94ZPpEe4Nic3rNdIwhL+S3YmkHFM3A
jXx9gBcZWj4Hq8f24VMlaFrFKXlp3sU22q1YK6prz+yCtatVdd5Ensxy0CM9wchpMVAIPVvpSsCq
kXhdIaiCwMcsOVDMFCKg0/E+lLj2RBclYvStxCkX02y6+8v1JWHK10Nzlv9e0CNDwlIjsh060VLh
hdfrit0hadEyKaEydr2BkF3+Nj+vsTlqh5x91j+4PA3l0GVvosfucJ4t6tNJvsUPNJvwuplFAlsn
Mp0udGfUygaoWIr1kXyeRkxvJVvWVlnZ02Yvtuj1pWoktyJQ9yw5v02HLysRZoiSWq4VfD0jJee6
8eYbQwPljFlcC0KDsUy1UGGSO/cSHaGhAQfQAoipUJGltbeu9VpVCqqHVvmG+xIF3rMrP4pw0Sds
UZq5tDYk42gq61nyYZnCxqH1Aano/5awOB5nvpSOM7NXfh+HQXgn9uz9C8aaNLTLSxiZVXXSeK1Y
BnuNV4QS8zmWAcQAX5TNxYirIzEIAkz/0fxsDZVcG2NnepLWdJMZLaFF8MDckStOvliSfvXbAWAu
PoeJN3cISsm7d0UJkPOiOjMQ0r85iWMStAuRgpYkQodps85Lbw5txXZ/BV/JpTgakU0YOfC/6WoG
tUdvQLyz5VskjQ6TEoAXZOA9DbdsKAbkb3tob1H14JBNH+BCiGlkDhBJLM4CUkuZPh6VirctxP5+
8KnGXVisThOYy0ksVP5NDUmxoZpklUxo+AD6R4QC0Pc/WzKvhX/Sl86L/neXS9qaz9pN5rFHuKSe
S0gFPSbyBUW+CuqL3NG2teSWRwzahYsAYwmWOJZccE9/IVdTuDoip+DQoPNf3pp7uIFbZPgD/2UN
/1aIh316BqY1wchUUxE6X3fuOIaGo8dlhf6SgCmtekS3iQ6h8l/q4XAdHdirDlmyH/XawE3V71pZ
a3GOVr044u4QHQJUGgYnhXUaZPzMHxfc1jw6aY31WAGIIgfcKmdTqQhb747ziJn5JVeGQ3137UOL
1Xtc4aSFU0PtFKiAgBstX+1hb2TI0WmAriVtjNkXbTAFXYo09icNDD8hZdfsCY/Rx7RqIojnIAdZ
fpl571qr0CZBUvpL6EPxAwmuXLKnEviKGs8YWHm5PGWrv+/BS+SFPZ8fBbdW7Rl5ONZRukWH9NRv
GP+ZlLF7kwdM8IOzfWjT3JfhVVdQ3DchCD4fjS8La0uajsWYyu+BLA2pIOcwz+hahf7SqBlzbzc0
3C1wPuV3Rrr9SmXWSEr6ukX6KG5Jmn1fTfymPXBfByCNpHuAZnfsODjElauostrXlWnkmEsAfB3t
59rCRmUqBEO+7XvHsoDWw6FABxODlSYZ579487eM9LL186lfIs8F1kDKu407S+5p2QfJgB+PCw0a
lY0zCIkADPnQ0Qk7sNf/avoFSAObdtrCppOKgjFh3LB+TcTp+NlegleQ/tlrKBvGzK2922QjwlIX
kV20oacboN6VcG4CzB/CWYRznjT4vrd+xQZpYSnu83t1I5lUrRm9kBaPpZIdddgwQozjlGa2kAKC
SM+UmxT/BrSWckPNrfnxXPt4CJaJi1JtHuKTVBd62H2JKnqO71GRA1BI+YIp8s7GwyczHW3xSgJ+
E/U56sqzU5x/HAQt3sYZCWvEHY8kMIuFbt9KVdCs7mTznMNJWGnXcDUc3BfTSzIu9p9rKLeItLR5
MycZyJ9EuZh3BPXeDjrhaRgt9qAsJNyXAR3xVN5JsElKs3BtoJ2cgxhtsVPDkQytJvt1UK4o7A5J
Uhl+XNku4/k+uEN318497f/DD05OO5h+0OjhcwLz+fOT4SvvtLDG2ayf9vXHc3OktcIDfJJodaGJ
AlxlASCXHRvf1Fhoz8jPyDhrrWUIDLcRbeW/2b1gfM6loksCQoysJfKDxU/yf2EUx7hOA5N6OjcP
wA8vn7AQPI4MAjFOSG4YVdUfQ8jvz47/rjqd51EeC1fJ5qsYTET5eozJudwHwgXpHH/dssftc4sv
52OEajWxHJ6RpZ5H1YCsSYo0Qj5s+JwpG33gMgnWRnZq6frFav89S9YERPtDnP3RdilpPVd5iH75
/8bH0BaedxqaRKSQkIWnsOLRzaz2yF4hwMYQD7qVdm58hobFa6HzPLjf08uboA21QRCWwNyGHUKM
9NMFsypbtLjbr0YhvvAm/V9t5DCj68qtNwXWyd+y93rKGvOAK5PFKFFRAZ/5ez1qkkQBm2J7pa+t
QPPp2EQKEilm79844M1L8ThxG72xcxb5XgG6tzNBswkPNGmL5HUPPF1+g8jJ0FjkQ15T0CRc5vND
NKaMuS18o9qobaPSYPXqWWfZr7pfyUYesiUSfGvnjD7YaZcPFC3v+dW9q0Vv6hDrVTVQucORBpQP
li/SKoxvIYpgcFnE5Z57vF8cDLnh5O9f7yyySfDKCd0rftdw2qVaTrKZ7KnFlXGYZBZ7w8ESsOqk
WSSLOtDuLmqhMvDVYF1XZxJGM+4b8S30JhY5+1y1bbv9UWWResRwKBWw0dk1dCo++tdKrwXK9sNu
AfGfuhxcCCPzk/D4tdWviG2E7Yg8jwyGISL0cyxGT9Cddqftuq2YpJgSukPVJ102xu2IWm6ErLkw
JoLNeylz1H1wK2KaBSc9Tpa3muofu6Yt4V0B6jpogu8lBVSZfFtnkGRXUH/Z27YgWzzwBgUQ5a+X
wsNuo835/Ez6+yhPsD4GWlJmfehs1eB56jLIS26OiP/cFg9FF0lHAf0KKWm5z1gHvwKMsSF0ADbK
S3U/NEJV3wbxEgD9e/pueurRrB+ytjUcgQSeRLuoF3Uno930OC2Thw98yyUWxu4SDSwNusC9Izt9
hekCXWudnviJyT7IfwJo3kNk8nETjut3WPX2SZYH2Kx1CUwWtbuIbWG90Kq2miCp5y/eGMnaMX2S
ju+5mj8t7OwJfLLh3IrAs3vrL7zjboxQREpHiX/FvJJWuCAomh/HZ+g5K3zUPqOIBQQyvE0akH2A
JWfbwTZNQOvkA8SYofia1KFIg0wSJOOn6Oz15OPx4ttjzWE4Z/aL9YKfQcUDycbhhPKBi5adGbJU
32LfwBV2lLRyi1Ur9dd+jrGuLC+aFvrUKHR6oXatYODda+LT1r+5O40ufcfK4aA2mqMkf/qoU9Ld
bMIXmzkZ0CqXTamJ7/ng3CRyX3YnAwKNY9VPHSKhrCm/b1P/EHxRN9DFlElVCZGOcnPbWTSbzCC7
8PsWtslQOSPGv9UCxVTD13bCju9JtQWN6yAotkGzQjvPEKla17NpKRU4O/OH1zh+lwaVOMKS2hfp
MLuqzd6cJTPylbafOqt0WBAezV3ZjQ5r+V+/4aJUm1Dd6Gl2rweNX6Or2B4XbySCOzhD358bogPt
kpcY8iPVzjtUXYdf/5y6UdAC549wVxicXQhMDgecnOmErWdJIjwX5Kh1Qqu0TWqQYbljZtwtlF5K
NvoTP0kA61auYCRPbbyVQXjzpy5NcbmbnKlBQS6DWsEyFVXGZwyepNrofQVehXNLu6cjZbIpjMcX
/pRpUjNcniN8rPbybUWB5AjfpaBBgq4gHogyK3/WoKt0+iN9XhaPcWY45u5f6KqvXRMIxtZEtcRq
W6Ace6h9YPYfWg+3mqRDohgz/M3du3hg3Cv3c6eTco1uXOUFYMlh7jpQcalR2kz7J4voSaH3fUvv
p6qFWz1dd5zXoY5B2CqWdzAQEjuis3RJfSj8uORqRPUKSo6kncU2JxMBwnlu1iuyfukWpPTl9sTo
SCwMCI+3O6avxzdZkbz3JmRtCRuL6Gb5RAF37FJe+wQDJn4KI5cr1kXsR4tBGdMbb7puIpuftL+X
CK8fntp2BweDEBnSd8eGEmBdvmSE+xYKNCnUfRC2x7z8dCpWXdmrG7nZYzDy4ddQmxhYYAaNFPys
MYgthPh7n2/1c/0xJ7vQ/+hij39bSPqXe7GT4VUyABYHadcZSWCbcyzVxPJ0N/FlZDkn6OmvGi+F
wieo6oQHExIlUYIx8ZlR0kDhj3uOZYMu0hbXFRnkZwjmZwkBW1c3OMad/muIvuyV32vMXI+1htvI
YZXBtrdVaukU0uOucxKb65fyLPENOJhAOjiR3Ij6eQsFwBlGQswZuEdjLFPIKCgQ8xCxytaMuY7G
TOLFgMLdQ4rnXboGKnSjj5W4l+zdrhUiIduz9HJhX/IRwCnNVb84SUK3pVatHVapvH10cHOm0EX8
b3Tj6bFW6D662LDQtL5xCkgYkMDLt1UsRHVQ2a+PgCeMrEIey5CLBVinfLoLSC5VJ7EW9rmB9A05
zYPtqrUO4qH0ZmlNF2J07ASIXeu3UzWCQnPaYfTN4s3r8aWuCb5cMe7eFMK0t+Hy2CVgdah7fm4R
lDCZZ5aB72pRZCyzXMveG4eOCcb0yRC11ejpnaCTulD9LHttXt10O43R4y7WxSZOUOCPAtDtGapt
WzfkCJYakCAjvd8ZYOMMyyHVKwDGxdH6Qe+xDzXokWmpL/jDHAZdyT6yXZFcCKegnTGyLkOLpS/e
k9jl6lRAWmSyThkzh1I0V2yIL6UJ3Ex0k6neqL2qblHtHjcV3+A1sh2OMre4ViW8uE+CjadLBnl2
n1GemZoSfLnMWu7GYYNpFwcErnKDfefPB3gH/jctrrIB9pzPwESf+LWNMbhoPyDknpyZTbD/NQLW
ht23XQ9vecrWYIQh8+73IR40b/B3hj7wAbVw4t3LDzjY9QJkQJTJLDgXIOPtd2MxtCemdaahEcFk
O4tPWUPDe8TjXEEicvSaRyvFF0CbIuICdXERoFcYHaH041npqVzrLdczf9Ral+IQjcXGJzIB2aGl
yFRj9Xhm4e6PCdmLMjSV6dn15B6y1/F7LdTHUNUhaM1JOTDRjwD4dsmH6avyJ28/eIR/+mzpbY6R
Jdg3BLT6BF9OXZGC287heuZHvfDIC+vcupt2k4lNgPCyjk02fnmkArQrjMnq76g75sofItx/sSqw
P4q0vdgm5IpWOgjLVetLutIqm4ykDlxv4TqENF2Uk2bFTmXen9rt7xYczljQAs0HTv6Nwm+aITZv
lw9/t06B1FIpoNckKyJloJdoD5Ww9LwWfJ1pfCZ6p+0pq06XpmWR92wsDH+1xvtPCvFSSNrYWKQ2
B+HYIlnXt/GTmdmUmQn5BGKI0VhJFIaDvZ2fPv6aklEM08Yg5MI6Lp4e/SJftjHxAoiYLvQdwOiO
k/aab1eFTGzGHo/wakTa/8LLDhKE5TflFypdxNXO6GeexmNZjq7K4Nr6uJOQ3vy0ic2U3Zn72tBY
W97eNdP2LYR+XMMVVuwgswIg9C7yhYoirYMLSjgTyXMhv0OuaKhZHQ+iH0UZ/YwpjfvWu6F5Wu4Q
oqs0UjlAqxr+e03ZdiJ6GQPq3s56fwp5k7vBjJFBkVhvXBLw3J+XzJzJTbuaipqq2XiykOq790Kh
6ynMqd8GYSrCwx4m1466Kv66iQGqbXYaCSTNh6+wC9bJ9WJLj3qFAncw8no3r6C+djgHnQEHvjOs
lsgCkTLKGeV1LGXYTn2vukGPhC3hwuHHLQImJqowh15cxW7IregueQvSsKAMvSd4TgkVP8MElOuo
aHSZ0Re6SqFDg27v2v9qbeJ3dbn3a7UYEvt19lGphGoE+xkKmXTA8gKDa+7UysNY4i9GXE1FTVJ7
wWR6rwyM+zTCMbEkLDEEkZZLy9vD18IImMSQFUhmiNdvHIL4ZzOF0dAjt2wnEEeg3OUuPGTLkYlE
DOHCc+n45Ys7lnR/ep94rTcIvvZCqLgaVqzAq7CJu7GxYkAVV834gDwCW/qIG/eaTUCtU/oVR52H
wkM3lEcKwm4g/peAxsC7IMZFQqRWwR2bUKkpc4ku903YJ/IDt9hIMmw5PKD5Rcj3kvEGyDV5taef
7W0KhkpEWqWnXGs4RxAzTw+2OYqKuLcYVI+3GEDWYk078eOCfFg+G7fHBsOh7+OtO2Nn6klgszLS
vbRJtz7eQ30Q4SxY9ci8dU77cBX6kEa0NbwasCEOc0QvFXblDy5WLU0kCho8/0wuaiskXGUdma31
F+lU/bj115RWI99DT2AdpMZyPemDohCiEl5/xXo1Jp5RXhgEtm88uAoHiCGs0H3aKhCD+i+IceO5
gxvnX+ggB5mhVfsR9rwk2BDj2NLjkZWo5LPnB3Q5DMvUtQjxEKZl0nVIi/GcBI54KQBFHFjVgwIm
aLgJ8yoeI2d9inATpZohVIsNDrPTv0aOnVI0V8btGmWEM96BK9PveXlWSpgsB100yPh/tOTuuue6
6IEp3QUsJPafOo+Tnx321k4mLWMVs5gEGEA59f9bIanibZ4e2nBN2UvzUttfSGrtlrotEqYOTGIk
2e45u0lavjW1XY4LGpR2yjXWSjmrtJsgViFgPDhFSsGLNdgLHTpKWw7Rv0MQSUz3SXcAl8AZ1kkJ
A1yzW2B/TxlyWPb2s/6nmAMXtrZWH7XS2cLnzbZXXHpwwwq2/WY1zSP6xAjgtQmFmPXob+/3kbKW
N+UaNffSN/R6AhPwQ3DqYx27VM8qSVn0T8olwOujyxlDVwfCZzGj4igjVvZECEdgK5Ol29Wd0kj0
IFfF9Knx7/zcoQ0wR7no1yVIWBfGGCA7UrNLlHuszo19aYwi3tX62B0j/fm4yhXjztVhBLd6mJHl
qLiirOuGt3jsZL+d/RtGNW+bFSR/mEQDGLtE6W5k9QOyVYfCvGkxx6LTxJHC4qdYTBDiZapCylcu
e0voxjmMOQuvxefMn4ess3cSu6dEPXfNRRheSwJo765qJTU1zA4zwGTsmZ0C6Wt74+yDjLgPkUDL
HHUl6HhjvPVpdeZuTIYW+hWNqFNSFdRwkHq+jKnCzv6WxupoWOlpvtE/npSs8QvNAGNCAiIHEknU
edXM0f0eM8Yc54Q0NyqxXlCqhTXy0BOGNn2TG0rBpl1Lyl+KMdfejiii4ifo0mBG1Bf3uyXZK0qR
VQcvEXeA5Yihm5KCCSmYX4CTDkR7bOEbj4YS/X7Lj1ELCfaO9RuZLmfw+aVG/KAJhsN2dd5tsZQ7
chbPWquo9PdDMfQh5LCksJCTseyFUdOP4xvkzUAz2YhPDHGmWwSF2wyJUF+XVsQMrqdn2Z1jmzb1
crpNEdmkKM9coKEPuvygF6IZzOP9WlSviRvHCOteTgftPprM0YFhX2VO7hODLBanp7cQz4mk+b6x
3t34fLselAS4Q52/WIIOfX4Sil6up1KYDJ4zTM5We+yOZkxdHNiVVhTNhi4EBqALQHR/fnvUY1Ub
4VXa8zsVFdnQ8JyWSj1lD5sNadmQVewDFyAHc8PEGpdFu0zVyo15iUS20EOkc0FIi1in/1LsVZAm
nKbcp7R+L2qOXQBmbXsQ1pfMazCchI4DcxYLNNuftsO37V7y18B8R7vdpSMvdLlnXZpZf8Y/sip9
UkP+w7vT0VvwFOmX1zfMwKuy11LwktcwfPRu7XAm/DEm5W7qEiZb9qgk1rM+wHlbZf18Uj82OtOi
D/2r3q9vxV7YWnNU7d12gGgRcQXvT/VeitrD5QM4edXXhEe79bxy5stsrvt5vojvUFNWt5tUX9aB
6i6CfXr1l2vVnWe8A7jeUzG8fLts9q5L4wQx5kP5wia54QgwaDq8VisIxdWVMmBZgDL1GBY5XfuD
jseQr17hiTHHxq1SFIlD7S61ZtwUnZBViJ+ShEP1bFAgEbmH0TzriGUK5u2zHT3Q1N09mL8naKTW
abq8KKNJNbyh+HB2zoUij2d954tE3WrxQ+JIQPzjApb8vrXz4ZD8C21Z5UNb0R/qFYuzRY/5+i8/
CY2bcVrfSwIpgSql72Ewe7wkbpSmgT/LdHV4dHYO2/C8LJdrQxx/Wsq3AEyfHZll218fhWDtdjpO
jzwrYdmwhUfiIBMY2rB7ZSxo0Lwq3/4YcOvSGferG23iR9+5UqvfBq6igfYsON3oLVlt5epzWh7B
nvu9OdRmlfyjMlg3FchqL8TI9NCL1tWhHLbshzYdWjEAdqYpt4EWDgeR3xub7hfc0dEZvucXEN+s
znDHwWjtveUk4ydClunKBYLr1vaXW0tCEv8xRCIpJEbxJN2HkRrgtlFqXBC7ttAfQa06fRbK8oik
uHuIRLO0ET0gzjiDpp0pCKmybvuLW7Gg9P64ABB/H2aJ8RgPHUSsnDPYma0/khb6hHSCFtf8ub5P
zfEke7u+yK4fnytQZM8ettd8ZhkeE9qKU14A/yUIOPQ8X5XVZgdPoVC2pc+TcU2087dJuOWTgH5Y
UtLdO5Cj0Mhnk1LGIlAjSpqwjTt0ePoGMkz/JHhTTuMzd425+wIetWA/MIs8ZCk4UkyzjtlUhD4p
Hj+tfRg/KcVaxXnkn87yFOkkpAsd+HizcholZZUc0Sn8VA5CjwbRgfmLcVW0d0yQCT7OsaCoqSB3
B2/1qIlfEcg+0hxbPyud84HoPDx6k8X9K79PYpV3Z0t/yXIDjtFa6gkAjB0eRN/Pj8gKaBwqYS8d
v3ElqXhA/ZhvrFiuG0iIlLcMgP/oNovza9FVWWGrBOec1zHMRM7zWOv3YwCYMOMnu+N+dYsasLlL
+Qho/P8WaEtuGA9SNClx8a6SAYcGU7wUEOfF7bqUEIHI33msGJ1ctGQty6a8YdCx0/W3cyyPb2CJ
0Abwl60gVzRf3ZWrGtJ5IRm5bYwnl5kQYBhjj9npp94vVhSlDVNly0hxgSwd34Pi7jg9rBIbZ0yU
zADke9g+xPS4XB8o/wkXWcFCNf5HzV1wBNT7m/5UmP1/r6YZ9BuLEeiDBssW1ciOFyB0MOg17ORu
ilV02WXCdT0xI8wE0l4610OkciF/zi5OjlphOvUqLggjLPzb5IYCuC02Ys3rnlRUTVsb7dzFnFjw
xXQXRjSnKN2RPM4YQx6ynJdITeYVL/msjCRiLfIu+OQViGWV3280F9APjpesSJQnyMHpbKVigq5u
QfWxkAQujxNj4AH32ks2ub8Y+ObgtJJ4oDt0B6RXbbY733XEeC0TgAHSJUl5iB9VHRbMfSQMjFN0
IrRCDpDJ/pm4F4SGMSmdJyP9kqlKlK4BgVbmCDA10gqTufRYGJSs5995qVAsjqnl3lXHiCPoVH7J
tCzEDXzwzoUsmpam/NxMlbH4pukWFAypUaTBtRKFkM6Z1Rp+2AWPeh/dw1gtaRJVyGwzU7SirzaO
ryvA7S9zqvVuDEq4+eGs68hXVgL76djePy0gqVwVvw7Cpv1HFpyAkym6hnyqyNrO8hrExTbp4/2D
lJ8eblvgtvYFWEwKUitZ3d1DZRgE3ZeondUpl+Ac5RCEJiU3A/Easzi0vjYDLkMJYxO7enx5zQQW
tBuLEuZ90Rm4Lsl38LqnbrdBEEZhIuAhxi2seCtAaqeLfWayB3ekfJVvCqmaosI9hK4R6lbBcCWz
Wcqc3Zpudx6bSb3sjW4LQrVj4K9rqbrFlf58PQTt6yPa5fx+iVFxD5NbYKu7E4QYYyms6G07iE5C
Pkk/hqpEvP20qh7T892M0kT63GQFDFez20uR00hmdodyw0/nibgO4qdqDCHCpZQASKPubN3aLjrG
FAKbYSWBGGd4mVnl0ajPLpNSFqn9+VkkhhlXWpR/GX/MsfDQD7uAO22LRQMIMueU1ZH/OtpiSUwb
Delrkhei87Ubq1rh+7EUr1sUofzugPCdke3AsxKAOIYKGBF3oeuD6xoeEmJxdQ6/rkNdTAtpLPqq
JzNdWSGN12llmgEcGuFjOs6ZSB2dtPXiTaAdA2ugzqae17IpK8A13o66Q4ZwOW3BOsvkmkq0Wl0t
DWmnwbxPjtMsfM+ccfZ18OI4ErfbWPBUu00MC0fzNO+8Jue0osCMwoIzmueOSwsIfeKxyjlU+ln/
tOPRJgpJc97/DsDOHf44GfgHJy26arw0F8rAVhAyeGO5DW8GdWcb8ZI0aD01Y0EnqA79DO1gXhlk
PhvvEwLdLrmXa9CwYnmGosoRCQyLPzgjZ3T1NfnTMiwUriyegrVuelLQ3TiHBkTWJixUIENIdrok
qSkxiR3U3H+JEPmOWnDldT8fX5EAyVL7Oi+JixLVQST+JM0R3B9J4YP9u9VEciUYrDAbvN80gFa/
eRYLFNmARZvFlFBU+5TvgGT4f2K/hfCu4B6zrPGLcsFJ2px75R3vsA00IrMLcTrgu/uUhSjTVUUq
LIPn/9ufvqz2b/TtjfqKWquNcePZo7FZNpAKPYVKXFzTECR/PqXGB6rdQAOg+M0s7Ayk89QtlvWQ
w1jTojH4x0fI3N6r+aFilvNUlwT76IrpKnC0u21aAMa1riZtUpREgwnSxxJLd3VqVtitWtwqeMUJ
ogmJBkSkA46Y9ZXIGgPe2TAYW/TWcsCPgRjrLzy1Yida2Ozz0eLOdOpepB/1wMVSl1ZX4BW+RdMY
HSKqlzZJYVc9tDp4FsnrDsy5aJNONsyZCY1eEr+Pn1piZ94qyhlbJirzh+lUBA1ogKe0/SAj3BgX
u3DJDNYbJmYnPk+iAKQuu2v0Y0liofjoY6tFAlNNNDska/dsK/9gkSh5kVgzWzUouubdZwuWi7Zw
jQ2FSICUnJOCrlzQbM/hpe/VjXNqtgu9h7TbYwVWcC/g7f9aNWpjn7BUnwcJa+nTaHReIBtovvv5
00dwkBMDD/Px8T+oxifMd1ymD8e7O/iJxTE1Ov19tV1NajHS0UD6oT3MrTV4uUou6k42VzX3oiZh
pxprhV8L+3IiAp6QRGS9P0qgk/J84qAs8iMBawHI9B5rjgYYFExs1MAPKbSw/tbMcg9fuDDijdNV
Yc9FMXbsVWH2cqfUIv2lTvtoZzHEj9//1bq1rEG+KGxAzcjf+LCU1WrmEPqdCjKSkwOaOtwU6kdd
bkGcAsfXUjuYMfCKeZNduUdyBM3w2zPwQrHfV7ZvlD2lOS0hQ7HSXKkNaX3MIJMt6yovqAb3LY8L
nIpgHK5XkwhfSHn/p9z50e6mUOOoDYEsZT5xzttdiCBM9856DxPMXuJjWwwqa9pxAjrBpeF1olqF
XgkT72mo/2M4aOKCQFpzRlmQrixiPHgbGepPYDjOA+LDW2rltG+mgc/C9+9Vr/1KtZRJLmvNbRAU
ipOPZjzem7c0QPCY6XyZRlAp/OzSkC0RKzlva8/tj1Hvy3n6jU0Zg+j8Hclrjvldn5i1mXSEgd/s
9kvpreeA8eCoMUEEot4i3JouwidShmblJCshJIeJOfOYLOncupWG/wkrvmy+DwvYxXvdx2rcJbeW
up0anVqbvUWv74y7Rv6y4p8qOFwlH15mQKvwB0tlB5QDSq3gHki84uJIn/LWS1D1nTd2C9+046Tu
ceMnULN/CyeDFL9nwoKJUsHEJsrHFt4ywyYVrKi7APLEn6OsMwH01307rwTubXHoOGx7dfbi4kXw
4Xij2ncjPiS8znblq8VmjODeghZRr5UUeJ4I5qLNgungvxGlDwU+B0aygChJ9OzDb7fBlfU1pnbo
9L0lUk/e0Efho+ABxzY6ZRWD/K9NXNambyqslxtPO8CJiLJjMgY9BfOY4KDAyCc4KmYBmgq2QdEF
JG0R0h+QEooj33Px/my+O8tDLyEiMTnWZe/0uOnS29wWG4wph03MluvC+YpQLiExat1WRlcgkV52
NTSQGhP7evR6dXRknIhyRYkys9GTNctpDtaDZypdI2cYCH8zgkdmOV8gh78hg4m2JGzhQ5rIL7Sv
e2vXJfAPPtLxKEu9mY0B2PH1TfY7Y57XRVyK5/1KPDXhE7dBkKy1TZfA9Qt9zeNR2rKB7DlwXFt1
ZA6gjF4C99G8ZPwz2dUbZg5Lesnqr6XV6vbOQhovsa3mBV01WKERhpI117GXbAw03jXGzecTu1Ys
EucFQcbZKw5mWKLqeFo2Yhspdl35Bh3XorBpfJoBBD5+1U0wL+vSyFkXabL1vhpPzB9FAipDsMOq
UlC35XLaIGdzV3vLtIJCnZ7FOiop7HMvygFiwq4takKkU+ouqeZrX9WdTBp7a/E/7LF7SivI0JhC
TfR/mab1d/NZL6eB05+HPR1jCDvhzaFojNp/SLEKzbDI4/1qqNadIyCRkhBbfmri+Ko9mB9YvFJl
B7uiwdfgxncguqGjAaTccqB9NylaaowDZfPocaPVRxt9bqSae4VSi7F76tLvwbQqJQKw8NWLonKU
CaMQhQKIA9WHJJAbWElMcUyaH5/+wJhYAeB1OopeVK2EL0eA8EOcPRY8yk5h9hD8HhVwSZkUwMAz
voKiuNszAAbJT9pMs85g87v8+tW+OpS2Q4v2b02tE7rD0nKNlrm2WW4qQQRCniq7Wfv7DLPgraDK
q48KiXWkF9WKYgk0KuYE1Y7BmzDo50B//f899U5kRlOm3PTm1RE/Pj8TI3MR9wClOKuzlQ9bjEcr
swBgp88Rcva5I8IH7AbgbQcuL5YTTUkDPCjsZW/32CU49qavjyWNGZvsYsNcZFFrTBOCsrxPQe1n
mGSzE8Vgp7wH1fPr2gPTcEkTKWdXm01DMSOQ2gWsmUtQzZU7MbnMw9Jihf0JsdEeRb6I5mfImPQg
S9JyzCuFAoybrGYwYz+14ltjdGdZocGpXmrJZ/yencbtXDYh2vqzUyaRF4utlpeO8NvqgxAER/iz
45qiJFawuuSSbBwn3lnFDn5PRhJOHNxyk1jF6la466blmC+WXkQSscI4CQ+TJfqvHu6mBCWZu/E7
DDVM6O4CpQO8d2qcUT8OjpcnNQB6dmwNxR/zNElHJ1Mwgw+X5hAqEQAxT/8ElISF0C04npOrILsk
HSeDmBFSE+EC3ZWAG5omyNnqJnWagaJBOmFAScQHa8sthgQmaFLgvVcA+oUCqdDHdT8hPpM64q1L
n0qHzF6AcJ7UyZmrR7e0WHFWp0fEbaNf9uE5KPZhoorx3UdrOb+DfgrzUKVwi6uJwuR3EygmN4np
ofdRAL7WISjFW5+jhLZwNNuKvnnkZY9AP0F0iVOiGB5tU8h4WvLXCxVc73OiwobQ9ea2m6DnWBiJ
QANEp6QGzO6wr7BtAxITcN5CBjLLZExVCN/zXMbCnRNpTbvffIjvWEENSWoH9jCDFiEUZXscMffw
PyXLqlWtZKOQrQ2sut3Or/4p11lps6EZdgiJdhz0OI/NGNT6vCzZPyZQKLIzIhVCtnaiNdNDTEWp
I2JX+sa73uyNgCu173VL1Dl2l9pDJXyl+n14IUXgVZ7kf5FxAtMjoh21MWBf1xdwtkCCk+biKt57
OQkxbqvCyES2A7PNiKh47NSLidKFOr/XroP0aKxljSQBOCe3uYj9UJCNgKJYDWSIIpf98z7DTjkj
YkEmUjaaJ4UffYGEdZsmdqI7XloAXjDGMQES1ziQoy6B1Bn1yQIcC+1dbyKXGYg6StXXz/hsFdKF
0x8AuNWvMoOjm4nhRTIizq3dQbcFoSl7XX2Ebzr5q3xio1Z/XtDkR67II8Zv4W93/va6UNMNz0Y0
JX/FQTDaIIBVD42UpZOvlIv4Vy05kIInbAwKilMR2JNqfdsRRikfcBP++2C0VQ52RyecSiKJW7zh
Nc/FMmeZ8d2/3ODiHOdmONjfo9XW1PwjGGrhbI4+wSUTlxqbHEyAv0Cr0Zd/PFYn+0t/lyyk83/h
JaS76b4z7BzBHmA+Ww2rvtE/4PbFk2al3Nx/jAb7F5jRYPW+3vD0NuGgeUGeZiNcYGC/LUMsZLo1
S4I8dkDcFLwgtV8dMhjCN1o3Q3rTX0aRNmv5nVP+0/syw7peHBd2+VFu35aszDMPe6Rei9YX/fbV
0owxtaUbqTu7jxWAPcskQKqquGxVHqqjHPDQgqH8RbZyFM7xcKz5/Zc7mG89vP9mc8+ppKkS+J9n
aQfOmdvbyIb6a2/zy62IW/vDXbH7UWh+4U+Zv8YU77k503r/V5dICxVqYndpN7QrUK4L6mchC5fd
HhaU9kHa1ORIZqqRbI6Ot27PRm1jYrFWaO3KN1jOFUhszysCoaYjS1782ZEXQIokqy66giD/6R4K
lR0OnHhhd78z0obAcsdJQI1jN5opoNJoz+9T6KRYaYH5eg93FcQ0ftHPQs5Ji9AxHEgJKEeMgXJG
oMDNBihyhr4Sbv8aeZzCQdyPgcnSbiXOdR8TaOIIWie5slvr4Mcps585Pg84RjMqXkXfChOpephK
42apK/FjnTySDuX+U57vHcISZa0fFKVgX1A9b0iy/sFudGfdpy8/KNu68yjcerZSCJx8ouvutfVV
AQskVotp+BSmJrqiG7y0FQAzicqs1iEzVMzQ2EOpyZRsT8DeT3VUIXYgQcgXo+0z4ljxeFMBSjr6
OTLJyNpW8EBEB5R0uwY72KKhZ9reHd4rFHZUnhbNdp5w0IE0FMgX32JB60E8h2R8tfB2CwhoW2Nk
ASyPTAd2ZUPewvnk1oQAkKUqyHIfUb3mezs/fyE8xpRIaotDfYCJeBVhfUhAf0WonQFHd9w29JlL
ijfmQmOXIqrVqa6xkl0Qp2JNS0r4TZU8wpb/IF9kLC/tsgCymy6O56jtUMEFaJhON5b5ZAOSPbB6
qKEyTJE5eGxy+gwZWJfxUZ6rGcH3+6y0fiCw/r/Ke3FB7d8uWVyQ5brxREpfRdPTmJhDJKmrEl0Y
MHQLetROcJIhTPXym+L6nXK/njsanLKFeT8diJv0et5rjUEKHThmF5vOkoYgRNY/m+CzldeTw3mj
2dMLiLDysKZv0zGZJGgCObUfmK950KTGAp7Eb6TTg3JlJKXCE15CH35QbimaEfw3ekAkKeG0egC7
2p776FS5y+mcU3oq7svjYzIwoiY20dFzD+z2GkeKnHAqYoFZfBKAiNHAG1C/3mYiUeVRxRvup49g
TDydN0WicHAZK5qXtoR6bsE//7YcN2f/K2McU6lNMAKVFM1fsYE4hnxaSLcAnNQcSrwFYfCdNH1O
ctM37M4jdhc7tlleTadE0HKBS5DcRWOigAv+6bDCEjrSKXQFVNDFMvQDhdj7sCh6eyRQTpg4m1sd
Dt0rbal2aGzuqHpZWng81AtXB+0eDxn4yfBXoiLVxv70TNCv/hNNyyMIyIJb8mo6XwuPCY+IHkYA
ubwBRTQbIkJQdfVNxq/7ULO/mzNb7jwtXRNgJ8vbltmreHj56jv0cQkzLuGuIOuPCQB74cV+C0PF
2Gsz1eZRTqbztS5jFwzv4oYRygmYtOM6GOyspAjUBP8Ujt6+2lf80RovVZOHqMOqgHkP2r9XzW2V
DexDgLncp3E9LXpl4h2S34QT5NUZ3/jDyw0Terru0fafEIpf8Y22Oa+BRc6lTSHDBbJU3JAWN7pe
Zla91JciCbkQjHqdh0Fj/aammtY0unhc8RsEQBXTZLSIXTDvQM+9JelZUg/Uf5sreMfnrgWZcXHW
PaZKDefkDpDu5s+p4N1epEzH8EyVyFpK5BbSceyDX/SosAQphXLgjuzYewCe3ZdKeBYgEo0ox9Pg
3N8ktmsHDPYJOlssMMM+VUN4jgUQ/7JCISJ5YyHe9KIL/tCaCJzx1cDuvOydtcrj7Eoo+cvTUEDp
Mgr+jrh+ksFC+mOrRMYPPeMCanZ/Qu7+FxEwa28zgycCAgkGNSaxIb8OzezakIuzC26QAiBZKWXn
Pyx9TH9dDCwQTLbdQc0//xGiXBUnbZkl7LNUKk732yvkXXbnuYsAC8bDyctegJCbqgK+Kv8s4Eet
/XBWjd8HFz6Fa8r+4U9zXbr1Irr1YksBnn4ZtzBQNzG2nqchTkb/DOe1F8wg9D+11HQYmVksFTDA
B9FkUA1RG2KmuipFvNEJnFI7Q8xpLQT3FrgD5EHIYPcjgIuKCxNjVKvPSROj+MKFgYKDI7QpQWZo
jpXeM89QDB45hEC74LhPxx0USia6epyWRrk8HnscHW7R/HVK+Ipo3lb+MGBBZK6cnicWKfvGuaJW
mpW3b0vulCrWRw7nwaSkamL9DvDQ2B258FY/geXAt7f2XZeqOK7eLmr01qCNOjjNLW/b0T2hnkNB
d4hc4s5L/EyFbeRG5ghZQZNg3xey0R3GwI4hmLYZFFZIVpUkfep7HgHNGtkDbyIatRvR3PLvPEZ+
iB4UB2c80F5vyLBKbpiOx7L7nxXBldTT7cSxtFcLeCxO+1kCEfrfspkGp7WBaxdIX0enaTaA7pTJ
Oh7YDLTG14UoECE6TTl1FZGG9cNNeC+1kitCP25VjRNlfqBQVuB6tcQU4ioCD0YxV/LrfzKjdF2S
gTxPYlHUNK8UC3BjkGz1Krc5G8Iyt6ldwkV4EhCYgz52j+ipG0uw8WtWtPKtPMc61ZyjD9c4ioDL
6KAT/T2KXmMkm/IvhnhYRVd3Ky+iM4rdCnj6Kju5/4fPE8FJ14xvhhDSzcq6C1duuYBN4W72WZvW
jW6EqHO6YOSnr/LfHlFPOFgmFUVRdWkYgrbzuLVypXp/wj2kXmQ17DC/ldAlGuYVxnz7FuO1A0NN
37fF2EEDV4jgIHg97ETWzJPnAs6PS9HS40iB099un+H04hF9PxErb+xj9Xc+lzPW3//caSv2F/Cx
DQ3TTwyC2dUH3otm8pGy6fxw1cWAEPUskUYtjTXEAQEoOfuALo7rZSnlXfeX81L0jJt6CsdHXx0F
Fc1xzyoiyUyvNFzeBTdHIncPtYHeBmCjb05m1+W46pkAfTSx9+s4wpUilQrS3fMkayhMyv/F6bds
piJeYzxF2NoZe03jSLtezV4fbJgnfqaQg+zBqogYGrPDGAV3hNOZY30MbLlOEWrjJ0XL8dIui6bw
ye41VJJxyBX9etv9+FXB7o4hJ9Sd+rGRtupuVX56+8aW310IHlnpIwbxre3l0h3diMepbIo4KijK
KTdO+tpHjZFKHBUFY9jvlZVOgRHLGmXa7VjRikDkZ2JK0ohvDVNkqSNq2/QS2XjfhI67+be4/KL7
JCrO6wc7hpnRYfa6SfFTAHAANN3ZyQqglNYppKqiqwyb4E1+/cyYIcQCk7Fac7Cpirt8YAJAJSlF
VKL4dC4vzdP/2BFp8Za5v8lyktJSup6pdhlFGGiWJXE4aef9WYPzqATHTgi16b2j4dKZbQa7d99a
Knxl5klGjp7thzExHjdyA0+T/M55uR+1Z5OiGYmsEDu2wDMVdrtQcTryinmVYO2DLEdNZz9g3y0h
TpSXT1Cw5h+pGHdusjgSy/mM/i4nJI9+J0Y1L+xE+fDZMZC1jDlwbfalNnbDFAIyjkggV2xesNDg
n9gUK90Jfk0MtTgTCSXS3+xi+LPrNmKn09tXypXtFbw39AeOMz5PeAWLEyYcuvkNUMyc5zVYJ9tR
tMPCn+XumGEv2vMw/9MjXiO/874IymIDSkZ1nu+4t9KOm3AD351jEnl67g6t9GhHY0q9yEwb/tUK
dg7jX+8tAfH7PZ6O/xeMe7n0Z1ghuU1c9DtPUWIw55bAtsPYUenT6AUvblK3e9VSUaziPKzXx/G1
yZwsZjOEsPfTiHbu4eg5vKOSyaBqBlaGR+e0ZtMiQxn2OjfhbNZZow+nowzx7VYZYR/KstT3zzmR
t/D9GiAInVIydXwFWTkIox8Q4RiaConNc4K7CqGjoYr71zCazupszsB9HNUvQ+E9a4L8+KPSKUvg
ESZzFhzWJXthNk1Fe6tnVcL+NqxwL54UYZ1HB3xsiiCWLRZRBrxmOZ4tst7+Llef2n+OFGEMUtFP
VZbOSIqhkhERJ8zc3NjOKte8ijLMIwN9E432tx/gaF5k6+y5JJjzqIA21pb9coANdlWC7hrhDqBk
QGPSSBErI3+qUE5q4dzEhjSqTQz136n9ZqcFjWT/IllGRRsXlcYyEcAlOY799RVwCMHEgNBmXZ/b
k2SV7TRcRgUsqAbYPkTy5fNeKq1CUqO00LajbuiM6vc0Z97/7ia0zmDLbvDU5PwNP7MwIT2HcxWi
o+mABH7LFD5oJI2zkYY7ZWw037+Ku1cKDWaxAdE1XpwJeriP3fGd93ziwAjqKtZufN/h9CNF8v5b
nCdzJViVx9ZENNBn3mjVMV4XWkWkWWl7HGb3U+t/U/Cevdjb8Klq43hq+xAV382KMtmXchyniBoS
k4CPcUYK1BFUqHbdyLNkIPsokq1FPq8lJfpGLSWSoHW8YVg56eAjtk/H8geREGCwr0YVNN3xu0h1
snKxNjgTUJlpw+355xtMWMAG40B3fHgIdkuRoDEEiUapyT5u1a80P9DsW5cfuisYVfaeUz0NvcXe
yAmCAd9GbtTXu9GlgVcyP17tLInU7RKvs1/C+sOLvJGOjX1uv+FdP4X1JGOQVSTtToJE+n4jnRt8
QCdHEVPr0xWu3vSmCWalMbwbxTnyj9Z6C3oAK36G92d9FBSQsKU6Kh2YMYd4SoGyPmy1mJDtOTKu
sL9E46/6w732DGQorqU2ucZgM5GhbvLRvDfCEUPPZm850ze5nlAW2lLtrmF60VktKHKtc8B8Dd8G
Ya1U0udLhbiTQbu9QRd/N8YUaEjzYPbPrQDYr0R9YY/NCFNW5FmZ0Gfm1Kh8Od41Iwmab6G5cSkW
6+/vxN40oUmzt9O1Mukfmvt9UWAW8/SNvTOgUlPbM2/YC+KsTse55D7rIHWbIE6x6KFqm1RbEsb6
XigpOEK6dKJA8uiEcw6SCg8RTbHH7gbkebLiMt6m2n/cSoQEkFsn/o7tKenjcj5x5jaipf9zPJ3l
8lmbtzabsJilyw5CMNSD00Shd6hPDjlrVl//fGQ62/THd+VZMOepFyJzI/QQs1sdH9p+E/GN4tOE
sH/qJkTaHP7of8rUvUjMgr/nH0Fj7C1jKj3Kkil/AhxeQyAva0mhtjNHAxvXXhl0UcjvV6/tVfKl
NguWXjHd3ZEmPtgBtujn4wIY2uWJw4LxAeq8JtymPO2hqHeLdj5MXD+RrntUpb+/b1l2QD7ZRZ1k
x6/5G9NW+YNdM4jHNBEoRCe09q8TMxzhTUCGVZzfugui2cW+5WftLzp4SfCC/OiI19zB0keSqEE7
e31Zs2kKt8RLWMb6M8aqeLRZ/nMfme4TXTF94wU6cZ4+YUIvhaEzqRcX0+ewg2wohiA1PEJ/uaTO
/LACHGk9JYPkXQpjySqGDjL1Ufjx+/DLFZaXp7sKNEbDxGGGF5KHeQZoLYF3GP9dp5bSZQZWHt+7
z2wpqnBsXrMolNN0ThPOS3RsNbi/82knQMcMrWlNfPpEfUGbBvLabcWWgDzHAJmbv+8L4CT9jTU1
OkyW5zFcQsCCS4TbB+VMsYiA0Ne8hhoRaunwAaeK2AKE3Y+MQ4KhpCN9YYIYidWi4b4v32qIjGEv
TDfPKVloAxGqyjNKZGD2v5pcOIoO7b/rAafGg8fz3xU8mADwhzcl0Qij/rr2jZkcZrbJW+WNJKjE
qpB93m09VpJBsgyk9B7mO50pLz3jrvlw4B0D7gc4XeXie3MD8nipQjrA/hWIhrdpfLfQT/MUEDR+
QdzGK9UDAdyoSYSZw4f4cM/As6WXcORLSv6H8zc77zJcNZ6VKklxiTVA1WsDG1MlIkZCOu7OD4uX
2ecbHeMAiJFksuxpuOropoI6PRfJxZVn+yp1r792LM4eW14yffPB66Lw9prrxCCKHgIYpPJcAsc8
AsOKF05idurfESI/t31CniT73Dz86K3ZGrug0NjvSr2ZgmfqyqKEFWbZA1f2kpKvxolr+U+hDbKF
HHwFlYxxXxsrJw42lyf7gFNcId8ifiq2kkKvZ8z4Uo9isw/WPdvtAMYO3KP5tRQhrjsgxYZSIANS
cGSwj1tai2XbniAemdERBFrVxN28uB7VuweLMlstJAZRVIc0evOcE9wl4ODUkFdsHH4qUGR+WhWx
dVHX61bczu8dYNRgrJoiNtUZvOlRqFrvrwwA8hv1my5kAxGZgT2FbkBEkkVc49QPNOCubudy7Pls
YuIBvepBPV32mswOktoGl443LxIvDUo3zfMxOZmUDApk5HqwrNjeImbapjFL0gAZv1FEG38h42+a
75dtfLUOnJwb35aC6CIGIge1WGnIvXUDubpwzejyCavVfB4kvCLzceSH120aGpGfqFOvY/l5aXBT
Zw1b/R2iQUT1lqJxmsydhQ5gLXPMO7gRYjvRs1ez7sJvUJM1Fa4N6I1kiRyHf7Euj8Ami5XIBLBq
VXlbz4/pozb6xoVsujKD2+ttUXtGQ5WYkF19A20SE4lIf9jl49i6KyaPoliZM/Wbue1ZyPjl34tI
sDQfVkkCflCfCJv6SWClZCxSH9aZD2kzXIO92X+bD9ku2Eei1VUT3Lc/fS89E8HoTEF2vvdyfUYE
MWHWD06PIy/0kwmxe2CjFwmNN472djXWKy6Ggx98fnEvoWSp8o4GZl7patEfhkoSSmAw7ryQnr1E
OGgwZihytlVcirIsd2UHZf1xLPvLYRh7fJdUkapVMSoipqkuGI5QOkyVYulITSD2IOyUB1wiL5yT
LoGjmc05qPSZS5aatkFGFjY2d3BgPZVUxS192Dl9R5V152BV3mLIagTf7JE5JmT1W9EUVGHjECCZ
PR+NnkPFCzK85hInF1nBziWezUnq+AQYmXbm8h8FnV2QLIursr85lPzm8SLULJPPqd8oYzXpxfuz
VAJBtSXJSsgIiS5LSxuv1XtkZGzF30reXKfDdbnOYfyvK0Nxz7u9NsoM+N4Ql/2twXSEPvvxc/xl
mMDCZQqU++nP4ELC/ErgCQRch8wlvaVjfQ4CUKg4LCpCG6QFLrM7CFEwk3ixNZYI4iH8zdOhrhcX
IxwseuHmQcBdPxeGmkn6No4JhnP9EEbaKqYzgzR3es+jwYwXpB/Q5G116agapCFXsFEjE+Zed75V
6PKZVHXa6hyT7vVpmK1paG3KrMpTEWpb0nFfhUcrStxVrIHxjkms1SIDhhiOmNRmInuHA+++dqGp
SKIXp+LxHTfvRU/mllcJ9lOW5L4l8o/EIyQd9fW0A1G89jAhzesdRMTsTdZc/tUN4eNxMsf8XWim
tzXxvi0g8cFzCQtPjwO22II0h1FE/pWpd1aRetcJVaPCYzd2rbtuv/aVCII7C+ImLg7MIA80uMoK
/ImkjyKWLSXqMbp7tEiKdE/IXRa+fixDNAGoYcb7KyMGmMFnOYgtJMK2AXJecr0aRaIE4eIcH2wj
R6ktJHCGd+a22vx0t6jBD6roMlrCGtJLnyx1snFy2H5JIG60lcdgAbdNOwDFTfIMEymolcvxjV4Z
Xr+piVwZhw0haadfdDkMFdzLa72vGbUcFe/3o5gB94X8ZqEVw7dfo2hy1rA9lCyQCUn/yjWX/rHY
f4FCekNVAJO/aslZ4N1q791Wc9JCzDAFp6hOfuLiVHv4gGQiAGGljrxhGV1oEdOn6uhsTUYs2+/H
sZBLnAv2kHmkrDb9bPE+kO+9S5gfP/MhzAr9pgrVquscAOgH7tb6YjbPNcJBVKsAPoiWl5p6ZDgR
digVQTHx6NhTIgX2kAH+vdEyCQu/wTyTKmy/OAoSdiCP8XK8iJID4AdvhRdTa0bmGuSHX/THUYc4
xy659mgt76v5LtKgLAyqfAd1fm/5cxhgOS7tJkgoR+5W23xQR9X3MyPxq6qvXGMrlsiErEzhaSvw
LAGY8gdGhYMBynH0JzQlamh92PMVqCnI9jq5YHzX6Jtf8DZ/VczCAyWmq9mzhO7KsbWpLhgX/VlH
UT3aTw1QCilIO6DcpomC9j8LUtzR4mIlSlNc27WjJAq+b1jBKijjhmgKOriNdieAk5Jq3PGUMgLY
AmOcp0/15KsaI/k6ycA/OzoajGbmLYdbZ1Kr690e4Bd8ZQ28WhpXeskVw7EplMZ+gVPQG7maaIso
hUAlq+19fE8QsAsO7cOulK2fna2JtjIQQ+4Ozr35xC50uNrxTgqlIW/X+KKcw5wJzyODNBRMAcCw
XAHcB4bkbn15M/9bKXy8+hAtsZXsqo53Nx4nhSYL+uxSsl+q46PDE61AY1efFQArE2MmV94shksz
aYk62vfp8wR2FE3gkBVvtH/5j+xhudN0sWNm34G89iUi937/9ZkQhS8oQy/SzsYKsPlOkODGk7xv
gLxBY+wXCGGZqZb32++83jt5iG1bP5zuvxelas8YvXJvcjB3B2GMmF/1WC11YEC5sLNrcvM+V1hc
qCVPSptAMaKEEBbtVU1F/9fYyFoZseruTBEPOtq1Co6OC0SDd+hwz8L7IsyR4Fy1qJhzFmDPL9vX
yV8kID0n1RvLxrCXMVyjYIggN2D32qgt1HqG9ZvKoCJq8e94K4bq8HK3/HsM/MY8OmGXq7HcPL+9
QMFNDJNWGqA1sTKasaFIfxug5yTYo5x+YP0T/iTwweiCgLu/yquocYWLwDeozj4GmULkWT7HOSsH
UYxHiUMDpKwm9HFpcROd9Xssw7DQIVPab/6FPXXY+5muHSrKkqUC7CklKo1VhovzD20UvXLWQybj
qLkGlCiQrYe+UCnbZ5N7iMCpzQOpMAp3hLtz7q1CAvTZzcQGZjh8pmoao3fpkBVmO2Wd8OxD+qUx
Qw0d6YHqFxGqZA3Sdj/FI7Rm/tVW/JMGa6qaL5af+LIQDR6rN+dtdDzrEc51aU6zem8dJoW3mIWq
tXwjKHSX3cPtGIji8FQMdELAmHk5ZcuUPqtg3kwyF8Fi9G+I3abCiyhI+z/Cuzc0q0kohf7jY4Wa
liX4FISTXn62sMssjNhUUhYBIhDQkNh/gI5bdvpcDOYWAOiBMVA4pAmqJbdWYaEhDgNl2+wSqS2W
7McGI0r6vqpQ9iaXm7uBK7RMoPGvXJjiGnc2QFOdWImfahhkSxNGOrXLEmVlj5GFZaLBeLUPLEPV
e7ZZIY3zeYi/3qtS86AUGB68iDT0usoUVUrohsQ0IR0H1Cpruo5qvK3t8QZ4UF1RZ+dJhN0F9qwl
CIJ/x3kh2GP4vZZUS114zX4YT5LmeExOS9CSqHf8EpI4KuB412SlD9ZOqZid0vxAO3QoYAv/zolT
6XDsyGGqO1aGF2aaKIJ9BinDPcrWRgR3gdFZBvcodGSZekxoAghcb36coSDfHZGvgVeJGI+1hOFu
TezZwTJs7+Irvv4fqAWrtClKu674uxvqyfMyFrksuzUBfRpAs691lqLx4gbkmLyLT63aIUYdlZ06
6zDAbDjK27GxbvQ0Z0uTbw6d6+G58zXaze1UIp42zhk1SGj7XA2/POjgiULIXfZckFaSy65wtJU1
6C08tgRv4LCsKaIQ600b81Nd8pNpuZbbHOIfUFjsUFJt/P6rX/aHUZlxGI6u/IFjx0K0bjlc7pTi
UsGkr6WRNvba0E2k8slSo0PAXMrhUPDWWPIod1byzvfxNC8lbSazxvuKxwWhBjUhrslRadq2bWgI
qCqIxk5SMSFfxfPz9HdYtKt512yokZDBq8LaOHBkKZ+3s2obNvQg5kxGjdReOVrHrczYQYwvD6Ze
mO7QK58QC/TXumD19+228wKfSJDnmBfy+xq1vPePpbxn2wC8BfZvkRxBFTCU5EJGJ4Q43E1aUcct
S3fbaitZlbBvdY+vR42pS2ugybDGx2cRKNjWJSiIxUzPn/mai76hxoK46c04qroGNfHgHwE2/C81
oB2gowkX+zyCHEVGQJnfNZfQcOswuWD8gj2KyjW3zsyBNTkPXbFAEXDuVQ+hPYshc5At811DZVMR
c7+lxOc8R6x3RZ1URfzK7TWZqwTzloB0sYQQuY9/Ttps22u4RH72fuByCouuqEUXKNBDmeO5qMKR
jfqTFCDI8qkF5VJegzecNNdioU/RwqH73xfOM2C4uLNt6qjB13CCDr31P++RwZnohXI/qwNMX8eS
V1LDbDtAaj/nEqxJqvqblGRBJyHBslOhEYsZA5ib0kjdIVHwaLVGjKWVIGVNzlP9DL+Ir2bT/PAm
lTqdtJ5zMwUEZSN6Z2T2lPmBQnK7XbnL6lK/v5nOzhMH4zIuUdKjJ2qh2Ua9s7F8fuKCIUzAYa1/
OXGQp4RD2jGYdbi1p17P3Ab3BscokH1i6PxePQyGNOUEEiYjHJIJYbOrLSoNUpGUyLKQGUvtdnwi
ZPLNt4TPXZGdNodS7wjpZeG+816QMjWJTwGHXpAkEjvs7u8/xF5YisA5LyerPVHnMAONK7pMfZtA
WQ9qq295nJCKFE3/4z630TOtGtNTpe4IAQ1WyUQicE4Y+GDU0UilSL9F8ZlfF1wU1ZofNTd6h/FE
E9oiqyw2wFvxQASTis3eBLy4RQXqFKIcwuyHoJbjNHFX4WMjTiOBRnV+cUVxJ3iTLIUoZ7KMTDio
U0ncqUtS0Ir7z9mrX4Nc6qDsdAZ3NcOc/bpxVQjzJYp4MhhIFiJOhyMYPgNPYWBn87io9f+euBZs
id77B4LEBgONcOTNprBGzUDMcIJUpNRRJnjoGSnpRnphnEazf+iDj7ch6cGaNVkz0N1c88J8FuZV
cjDdPeMjdfXuu8sB6XYb6KzpN+I0JdId6z5di+SIu27dpDy5ZctIJKAXkPCHfHDvP0ND9wNyqHVP
8e4F9pEvDKdvYYv+PF1cHzuRLT6UqUvj7Vmpc7gdorPof6Xw5tgHcmVYB8+n5vvS81hXXpNQ4UPo
onFcRozSQd/LgX95AfAh4UUh0Rymv+cUsYgfwHkmbjNCnWNVW2DdjRra4o7VGugFLq52df0uQQ9h
FaiaoqQL2pL0KuPAkvqciS8SGjiPhN99pJzIgUMVv7NIc7uQTd/Mw+/FNUTXshDRmUSJ7Vz0KuQb
9W/sZ00aN1YsVG9ofpwPISixDk+wTqIZ0kpnUpVgUkVkPBXcRNDYMAZjF4sMDSp5/p7z2jikM6C+
vLxlzFGeStno5UwgzcdWLWtwjcuvYPFxMDb5nbZ8QMdLZsdbO2ynhQpiMlEWwHG9cLpQ4SjYnhV+
KJk+1mOuFYzOOiLen7y7NDUc6lSZn2zpZW6cdMBSHo5cIkGM7dkZqIGzTTimUnwjCrxICSpu2Mb4
qprx9qQjj/e9U4zORNMNx36DInLZqI6qAaDubIRHBrYPReJ98AIjaI3PscEZHwLhkwcoC89xHB6S
IH2WZFQGBCDN9TN2O/Kw2l0imQpuZGSmIjdif9jurT8/Kid0mw85E8frrkAhyOKhyqheKH9V7LQE
PJRVC2juO+TbiC/v4wB/ikZF5rxJc342vO7Y1djSMle5Nkcm5GQQ9+Aiti5RRe5op/npc4brWuT8
Lf+YpVDZCAt+6v1TxyOfgpTZwI87L0828Xz0YX0ooSqjxY73cxigqUzrUUFNo1DZef8vdDRwb1Jp
7PgB3ddORqny6gNTiZSJ29w/wSqPljkvavj3Pqmex7+6oziEQGc4ka8CljTdpn+3hrHTvQD3PcRE
mGjWnDIPmtEZS+lM0Ztu3UQnpmq7zSdvnKbZF9i9mY891jo+abhtOxnlq59E4NZE/UXsX1z/EPOc
SNeZcD+DI7N8cwDLQkcDBdf1QO0TycufwLe3iqRJCy163n5SQKzFbiqT/HsnDzeg//VfCHq2zyFA
yUiQCiIaDOAQXTdRLPjJGd0QO51D7IKFewNJnF7AgQvP2pfsLzp5bMRkH166nmVWwgkeXOCDk/30
oCcHz68Si9/B/vS7aLWphPHGvg2n0QMUwlStaQil6E3w5ThlkyTBIi1o5CxfvL5m8WenGkjyPd5w
KMb+tlWvgkKVdZYda6zcS7MeHBOhyQ+H3xvofQkrNAx9O2YjvHiONpwIAqvbxY2X7ameW2PTFcBa
bP2moIMtvBqjuUGLMpoUhjp8g0xgoFalpq+086wNY4gonYq6Dz5fr6VlNrwSYWQ485jH5Bv3oZ0N
ezaU+Gc6JX1kGSSFtfHvrabHZjPXPj9IJz25vnKVgOM/NnYjCkHHxGSWJCl0iYCICN6MuGYmFalQ
G38aw+/lzBx8XiimywPULUvgLXEdfcqtsoI8h7LQqJOUPC6CEztIWjAWcAPNgqky+/Q3b1TeFan6
A0WDqhn77AsRiF3YlSMLwh/h+NKzitbWPBFrHWSq95nkkx4OI6rJMOphNlGuZOrtCT46movEPZeQ
szwMNAWUngbiAsCTFqXVi6dyIjgmLS+vxxb357f7WPp3+I+Z9vfO2NvlGrmICDCDikJNn3DFez0D
uQle24BN7NHLrnkKnDFkhFPDr245qXrEsJzHZvXC4gOeSavzJ+5Das0GNNgoYJVXGzDlhfJ5fNqi
HPe+nnKDSr8S9mGUe4AoUQaYSXypHCkCmlYttmZ5RW9Tj1b9YsXX6WmKMOB9ohYEZdfS2NwQuaSC
B6S+mo/KwbvL9YMMdpd0d1tK5jrxyzmhaxOwMpMHYCmaNykPw2p/QuWoy/GL9HQn8e3kNr8wlxPB
GhC53o6w5WFkF8+PwS5iqQW0KMx1mI+729Phm8M5NCzrW9WvMaPwG1CRu58rcworhhisAeMibmW/
LigsFLynljGu08+ow0jGepCBrwtwvMblTgPnF3HjIOgT4xhA3JF+K9Lk5JbU4OKObo4E9sqMyAb7
IO8ODmGtFmHJE2J6aPQJjYExP1maZbzwOIiIcfdLvWDpAbpQEh6m7PWf/bTUvawX4+AZg0ucmjLT
2/lwpRrJ/mSWVOl930iQnP4eVTnrW6dNEeZmddytpBTRX17zOPDCMJhk9BdjmfzW4wWVv5AFGFPu
mzIbfSDHl+Tn8LPZqv5rZNeG6KnoPJ3l6AUayU+3K6kRoobqTMDHpDMhYdQ7BSmZgRPnZyweJs1B
xRFSSPy1Fvw3NdjXn8St9ZHg5UwXDE7CyltM3GqS4TZ070uJispw6A2aAgCv4lpwQcGTvBTvKPQ+
dAiT5NRUNJ/DYhejvILtdRAhImwOCb95hti/KVCGoL3Ge1riziW68Z75me1BgPBGybfAJNS17TP4
vNr0riQfiHZXolSiYON+IeNlTlvwE3PmkZlc5DRPlqxZoKIT+7T78t7gvYnFnyAh4o4LIWrKId9h
7PickblxcvnElHGjSCV/EIAlQToA7QVEsaVoldN1FQKQ4De9UNv/H6C7R394DvJA4EWN5aqJyQVu
okj+gzW1mHINkZdOMDSfo/OswDaX58DrbZGz+OaasQAhczSrdcfZW2S0MMXVkFlXsYJ5egtHW4tS
5sNnZzOvquLkL9LyKKTq5KloIF74qzlbsn2hzlRRMSHy+h78M5070f7pLUc8EejTHbcZkV679XTY
Eswu5J9gvuzd4Rim6w3enN+nZzjL7xywoLgEZHNkdI+5UlPvlUCYV4JX0Cm7C9hyc7+5cyodzCqP
DQG3PzpvvrAHgLmVfCJS99yY6heks3fkmjf3BSffLQO1RWVFCvfVkTuZkmIqjZaiM3P7erlrMRSL
vvLcob+FzTG2Wrzi400XbBTWXVybFfOLViatQQml3sTo7mO9aAkArwC1uL4JDJwUa35nb6r8Ronz
fxA0VDAsILRzNAA1B9yjHIlAgUu/BdtW+PrCR3aQ1LefNnINW/E75hvMBKTdm6eyFRuGgViDMdtO
PLdfnQ1xZktvSf2jk6yHA5XMKGn/NVPcpB6uRs38lkoMSUFcmsMR/0ISqYxb5gTUEdB8XG8x84dx
VA9GMectTAg3Ypm3il8oiLQCAcmpLYk+0TNYw/Jddla0JHEyOQLHlBKDo+GbNeLldVFcq036O3Ij
ZV8BNlbQAhKmq2lhgh2ZiZDXkmp6CwC/e3Cd/3U8nBKsSsvf5WMLQbXNRE9XI29f0YRwkzfiRT3C
6uf7hpHQUUayKpLukm26Gw6dPy/YjUpaN2SsmbXuJXTY9xZkU4jLWrgwCag5BVz33jtpLXXbhpCJ
HyAR1rcoZPlatA66hmT2aFuZ70LH08dE2sGPpJX3aVgjufTdm7y4ZWu5kWm06yurcLTdlcWgvoDX
mrAWuGbRJBN/d2nyKRAncC9OG3k22qXJbaKs9fNu4tUUnDCGZbiuVa0vGolDEvAxUqkN3C4MEnCi
CqORQkE3zNZBcnG474vyl5ivrs1bkghS+cTIo4FbZ+FKikvj2SF1bzdZwj05IDpsCKDxmTX1qKdp
BEiAr+0kEYdmf9cXP3tZd6zkVce6UQIJIo+sHv2bfwJCZ/VK88FWlguAaxoE7r9RBw3L+htFnk6n
yqj8U+YyCbP1dagmebUFYLwan27t9ALFJSN4sya3NZoOKPVKpTZndvQzEKQM9QeG57Sr2bPFIbaM
pWJkj4nqR2xvlTu5KTgeI/SOd19NUzxjZ5q4t86Y9EFP6adhPgxD4Cu9Si9S68Yg8e2zbV4hxuly
ozjfR7lI0JbnOsp3PCQa34MGI6p1KJaeKV/nvx0jHtfck2pUypvX+GpMfhfUaPVszfG8BUsw3nT/
oSZcJKInB5vV11xT4ZhSEtLfjSxSU5wvl9SBhySVcUF4D5FfRDlH4PbcqmjKBtTEo9MfV96uW1Ee
3dHxYuMrpRw1EB2QlWJeCx0tT3U5GNAnbwaprmNkNy88tmfdP3oXWiDVgElfNUcK0em0md1joUcE
I9QbdL0y/rJEqI1HJ+U53zQ3ItGHqcLrPxaL8iHqu1mm3uMBfzrOgtsrB0f+AXCHa86FsX9UwThU
7Zb9GzohWiseSxL+z8mW/aozdjClZA41QJiSh2gx9xv/H3vCjxFaAeQ8uC5GEr+DxF8KflQDSwYF
d8XsWD/KMzE9NOhPleDKENKfpj4W1gebUt50BXjdt0q14hOs/isESYAmZRoEWC8O9AnSSMbH0VKI
+2M36Pe+T/NG0Spux1Av3HJe+f+RuyyEUnDz0Uul975qmqzzw+UJPgLzSARAuTouPYhXoCNnS3Vz
aI3MYXtLqf6yx8+yn9xk0JLXGHZI0ntYUJSzpl0CeiEt/ZVfEp+2E2uhyyywSvx4Kf062uGcdCgI
/Y0GZSvasgj57U0byF8qN8Im2Q4cW5FBCy4dKEy2u7E9VP+HLX9JtsyNntUu37dOCNRSlmDXe39B
3/4v1XvzMNrne3S8yZw+BjZGPLScCTimtMsifSofrBLTOqJ9dME+YhuZNLiPiFPjvt4oR98gJzgx
FNd3uP440oMmJHhPr2MwKJi2HyBSSxZRBLw6REnirKfTZgJemJILLSZBB4TOx7vbJwK1WAzO2vdd
gK4gsqk+P8q6cUbeb3XypAQ5aGnGWuO0KYj07SX4jSvyH3wWlDPGqx0/LSOFB8wRgafxPjqJa6Ym
OyEgLMNlFc8vKLAEal7Lj1R23VL//r5rWLmYmnJ0r5js4e7jjRbLD6Lcrs7302LOYomse5A/xZXk
NY+DrJfAoMzQRQ1GfvvEAqlGKaXtby8zprcFbdkoEhow/TBXl1XZbtmYwA9smmclaFaC86pvT8Y1
fHdIUgYGNH25iOwbt7FGP5yzVv6s/VcRp/tebf33JY6zPtzdjcUhwVN5NNbWtPhctXQhIa3fTccA
SE+JaDljVz0N4RMCb5gncC/NCvEUixhPzCdaD5b1JDn6zHDOoj0r6ozTy6ODdjFCTPqDwYNZ6hhX
DpnQwWlVeu2JknGJJDmY9yw1wahKmkI8ACrCnVmVNtdoJgo1CSSaBRaA+17FcHJeZ/Ku/xNqeRzu
0U5EjL7piY5N41R3ln11ZG8RmHKU2z77WFICtz/OazKMC1E9WYnOFDm11IyTHvIMDkutlHvyJx+4
TPoNPeQPVLHOFSDGEKWDsAuLz6GhraqaQU1gTJJDSrEFi2XB4WssC9kkFet1fIS/SscFV7YlTTp/
/AlfM1/DCcA/POJzJ5wCh1k0FO/Pl3eKIr98Rc6jxJliLb9p6OPfTkFWJBVA9CuGRDhWrfZ/1MyX
iwFClbYJaJRTFuTrVsGHXKz7ke8mH/BHzTQGTNPHAXoAQND14Rs2czg0x6RB1KxsPppsvZfmK/v3
plFUd9C+tvYlFAgBGaeYemChfoy1K86m+MVLCunDvkCLjpsh6HOed4yVHLcW5ifmpMB5G/gL7o/b
8n7DcvZNgPIiuh+ikZv/RBsTsA6dyaMFqOhUOQk0jit1ddwne6+oqBJ2aXLWM/YTt6Iu3Ct+cSTv
8Ukj+GCXdawVjEv9sDr/KiIwATO2empCmsyifzJKzNaBfGxy5vEc5jn3EJkHqQzOd+KJbDHt/Tzu
wquLoBn7uxa/m3vK78EEuLCJA97eBjJ9avj15RmtvgtcX0pawc+FBVqQt+Yj0Wgpz6Rq8t3TbVv/
FpSEkcUhFGBjTyIrZvHH3/zlkMWTT5GkuU6tnNu1B5amCD1SsY5LYh3GoD7kBh/4xkdOryJSwTYF
cQapJvw13AykHAA50qSfNHsbwPVo4jL1Pc2sDHrrmGNigpw4iUg2fjTApY3NPOC75z5ECnbhgYfP
iDfTS9LemIRHoqr6pdgYimloCBr9bhI1iy/p5RrgZs+kONPeDhX/zoTibpxhb1oeJYlXAZuuWmsU
ySp9Q/0hwXA3rc9ws85L4yyUIpQuta84VOrmuRmlBcQU5qwiQtC3zbFES/DV5CL1f/eni3RiPcXC
iphz3jA0OBD73rbs0OwbyHwhxBoSKQI9kza4jS1iKKBd7bO20zT4dsajTXBVfbN2jsrmfkXLvU/p
kPMuO4LRWFOswhetZgHohYKTTpo0Yiov5Xg3xcafOtAJedwoYyw5TmY+f8keKnsDLQdefjMITkiN
QtqSBBTmEBLPsExFY4cbvIAwx6TTakZv7zYdUo0a+qNSg4jiMhua/MbBF0qckGd0E1UJXP1PwcAI
e94uhBVjZajc/AywkXvaHnyFf9pyjRcD6sTCwKpYOAs6mFpnh+wYjHsqzqRhk3ApUzW8IYwYV2oM
SzHWob2W5bGeJRzRq4w1iR1Mv+bdy09EFoy5+JiJ7X/hfdpjVm9GlsrVMmWfAlUMYZvyHSCUlG+p
RVkpbzCjlzSdpdjs3mk+7HnYoj234McBGJ6Fa4pOf2LPIfoNV5AG3FFMB6NxbZZip82euj0MYQIe
g38oOdIt3JCBnANhHLr41I2ROLg7MFieBjiuopAnqMeYxj1t65Vh7jqhlusaWuQMrVfCGM4Rzi9k
Y8ubXNcjUGrp1lzVBq+3Im8sP/jHkOAIwU7k40IKFwinYe6Tt9XqDmlOdAy8M6c7X541gRRTfU5s
EXh16cEBanQcslbe9DJbR35TKUBtO91IPtoB6bQz8KeAam+RqVWC7nX5in05XiVNun5xllh1Pcxy
sNolmxxZp62N025dwIP6FijMbaIOPB6fHX8NSfUoqg/+RUbGC/n4RrjxMh5C+2PVplLZdePchvxs
SvinMya5/RHCuOJpt9btcdfqjtmG7LrfrJiim72S3nCI4dp400DHwa68l6StrHFE/EwS1xzAXBZn
NyjBSMwbc/wsPllDu3SBGgE0CLenG9RDrG0i/edhuO7XR81/B6tE0DQb39sCtCUXP0EorocqaXrH
g6xTIbsZ2zosj8KxnWkBB3qoDZYhxkM9cDJrpNdyVz7syXwgjISaEQ/FLX9R9LChSnLVeHsheQvM
0grtmOnKHgl6w3CXfmgqqL7sxhsfO8hUTDvTayY+b3/R7lLXxB/2v6GVyQJE3dbT72aRr5oVX2Ea
0LoHwKzxzd1fgLGnKKY47bdhvoicPpmUWAPEpxmhRLxfKEI1mr293+mKZ7ZTtPAgyP2iCSaKNfKT
IkuhgcjYLqyJff6OMnJ/CigfHSoUvLq2f9WjKl5s1Od8K94gaHsUMYpZglrmfxYPlxXmZysa+5VO
SLnzYNSvyz0S/oj4dt3t17zutm+7DJcC95aPFWcj/fwQX5SQB1Yz0KC9N7odU5jE9luECNKig492
WOpijvYFjNOfnqniWPjAPD926maGWNirMFrNDGcxNTwmJUvAB/x06T+Mz0M4lfRp+7luAlYEwlsq
BWOqxwtsaRTNfRdBCoyhVLhIaz2r/S2MJGle2qRiWVaIeV7623P3/sGRkUzSkrWExgPyAyna1wue
hVBE4Ylx8fw9RJDEnsKVPc0L0kBXlYy+JOfB0Ov0blPzGs7jfD1zhDk5SoBzYiYzISDN9UxbPumi
fbknOI3ADwiz/UQxjg3I+KISy0n6t7Ve11TjengrMHZ04EtIASlK8/Wx+nL2Qw23NKMRKzdi0xmq
M+i+QhWU7+/UQ9HT2U5KuXJBiSwqusl2bca4jFfwBeCQHO9qOSnkBp6/gT2AT8ZJcQ8oCB4IG2VQ
syNr53nn5UDmVAS7s2ZEXPHd8cHcnnZGXPBuMRoRO9U0fzlDoGi0mFvwTqp2NhHLtduixw+K6m9R
69C4U73sxGB/dYhlyqIa/fEPuIm3bROhwxLIgmlI0E232qdKYrqjWeYpQW2jW+Yc7x0HOtzEByL0
YXGBA9/VAc0OBPFyAW6GvkH25OKIm/3VknL2tEldg0M0TwnfVRMqF+JcUKJol/0tG4kpXhtsiPqx
1+u2WiuFEOxJlfPKJ0zXhnJYJxmKmbeixDp5jVivwK6MOC6CffBIfXJ1Yk1oPoKWO5LwElg8S0n/
pf7WNup58qXalpEBZ4AMUyFY
`protect end_protected
