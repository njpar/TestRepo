`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Do1rO2c5wPIkTDsOW7OLHLo4j6YzfTkKqkEKT1nNoZ4SKZMwxTOA1ag4di3GqyWAxndbgQdQ03KR
xvvYfSME6w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lrS7YE05ZR4qGM490L/rpbUZV5st6Aj1ehu3Yv6Su6pEjwzAzM4Ll1KY223UxCNUJOuB1Gk8C2va
4kkhP9QeslS7hltcGZVkE8MCnif68mPbOPImaTgGNxzoof6hZ99Ktmj6wMsTqzNhFrtQ9e5bKnBo
YnFqbJ4PhKuBMw/ltxY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ca1TtQ6/884P9m3D5eRKTeE064Nd6EUU0pFpIqodrqHkHCrOvUvQHsoUPAurFiuYcqd5vkAq//zU
QadZMfMkWANIShylDLuMuF5EQBP4ojuKzBM5ePXa3di2aBW95bN5TZBLdZupEM6WMCXqL1y6P6lA
oZkmFmMQOOe5nLj5Hk8SvhaVA7DbN+qhts8S8n+hr87BFjzm8khszKAixA2623ulONYHYxuQG9rY
0I8QgXqqztuMa1AylcbY3vPn7OGr9G6YSEWXs56RAq6Ku6wNj8Phli5ylCsT/5XohdLSqMFG1Qx+
NKiV2njxdZUK2CayKQpLCPqcT3WhFuNi8xOTsg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P07S7qXU0u6S3tw55IySe1oMFh9wTBH+oHfwjy6BbJORPiiDQjMqw1cREwxtFCBA4BvBnpMCNO8r
Z2cVwCrNXVYJmHAZFnXpeyJcN503tZwshNoYmAugdoQk4JTfNw8qx//+/JGecFBrTtxK2/vaBQ40
W3T2iA95br/1E1aXp7oCt3ej4aDxL2pgJnEzO4wfLFfFW4vhIUnZT6xVa1kO8T8JsPOIyVxLyAh+
IT3xJRaNiuyYSeivKKMMrwc+Hm2SPDmuwS4iTg5tEBQxiOb29x0nYCHUd0l9D6zZ3oVZppTSFERC
3yt13kIT9DHso3JMLKChiEqPlMjLvxX41FXo4g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ij8aWT2KAsI9E4dMvJpG6GdTGv+wUF+YbVXm8oDr3aJKfSOj7DYlqMH89T6p2lIdOLVMiREWKh4J
Xo475NGlrD9PZGTE3cPgnR2IqLZKe952fC7Cc81FLBsc+CSI5RyOKbCifkY9i/8uLAnCZ4es0rdU
kUrP1029v0vCSFv4ZG3pEiEIQV1m0JKRrU3jANW54l6AIGFPZTMVtX9/6olHHzHn0oLjWWhYjoCk
3os7QWOKkcqxC9zkWtnSOgqcnIFyi1M3vSgrKhWhIXVQkfHBpMqXX68aahLwEU1hv21Ry5cYbPb7
QAxLi8ZHPi3ZkxBVg3CdxFp5gZneE2PSxOLxfQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oxyZvTqQr9uqmwIR6iNkne9JP9bmJNM6cn/MvjtyXri+EFftL9Ieyx2s2/Lzac+Homl/BRNcBBYl
1dKGt+g5osq/5XNCfmVYB8I35YM1s+kVSkw2TLaVzZ8DVkw6Zp7qTXc4szTU+Q+f1sKdvoTMa8YA
YsAOx0UfXenrgnaaWJE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yp7Mi7u4sYLm/InEfyle30/Ffcm0UkNDR7EdKiLwwxttwbJesAlS3rSOmV9BePLyOLqHLf0/DooB
baT6gVWiu5UHSF3wSFGKnjkdY7AUTGk7XPJSv9afer569FYIP6gIMc+LTm96oEUZYpobfvElC2ik
pqqVAfg07wsy49XwsSAzb3MwIXZnmcaqKCIws5vI0pmbs8OxtPyXRenyC7qhK8FYLWO1Ong0wecj
Blk9GgWZfKjkwDrpo87YOvOsTzKPdZcMNUr8t10nHDYAi3mkTUruUPnctXOZmex5jEtY8zxWWl2i
mdiXc5bF0IjD6K/wINDE3PzCMqJO5e/tNUhUyA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 134944)
`protect data_block
dY7BRYi9NGjs0QGeKUedPr35i87g3e8LCePzcLsqeXGMfPiLhCqfPGw1kiLKb3jCh3LalEqwoznC
mPn9tEdy+EF6PhoERyD71kxD+7DH0lZYOJ3gQkYg5XdcUDGuONlSRqVRjQZ1PV1zYxCcxAPzPpFn
mwdCL88QmCnfG97tZbFC7rLlWpHCVxPhrUWjmgCavtlablFbAn8k7hCDJKxmOzwW73us5aTURVby
UhJyplqJOTc7TThdwghH8Tflro6/Af6Av6xdZxkQPHd+wZ0HQCF6GlFIFECmfqp0Qf+NpMp3bO4e
cfOJLLOhfxpndtIoktYSh0iUQiaVAx/iOUUdN3e2WNbVzJEGzGmwRv7WSXgy5ZA2v2Pq2ikvgGCb
BvYl/J4d0DI7LyxrYamJ9uRz6USSzX6cUyg/zbdHykXxIphmca1uxjf3bUlbl8Fo850H9w/JiVtt
0/O4gTHtTL46QP3W/p2oK9sETQn5E0IRAA3j+449R3ABlEVvDMuK7JShCJDIr/WlYdbh9bgFATph
G0v0Efi4LoUTc0j14LfUzNPrnKgOLAOkyIbSWaTdEHZT/aoWrfRiHE3Lu1YxRDpbZxzl9EBO1S+s
BnRwiWQGzor7PAI2iVK4uIL6g/uxH6sr/aksCObUwSEs3xhMyvOvwaZFgw/cZar7SZ5vACXTJeci
S4ORpEipiNQZxlQyrvqYOSRRYIgcw5VsnK98Te4tPiqJJlTtl8ffOwgH9Iv6mld1+kyAVfj9U7o8
aBqud+PW+H/um+lAkeHQjUGbyAS0k65fbghjUBVWP4w58iO/4HzHd2UXQ6IvUhc1lbGdUZ636RDK
Kj69lWCJUs9EkZ325g21zSc6OhRozySd4iFKiMvTLrLhbJhXeRW1/BGT3L7CSGzaUMD5U/anJTn8
cs58vlOOtV/DqGo7UFpWZn9487dD/SWIjnNDTBuMWTtCKGyJU2NlE5YKgp0T9UqGflc5IOZwkLwf
71TFe5yV0roA7KWYec7+fBvoOvjO5BIGowafXh2ULETB/1EYOJ4HSqQKnoWxLH9WNObpqEtf/Sjw
NOtS05jd8tjnK1qWGuDJT/O3zC3E9m1vQJX8hZeHlUcm/9ZxHwhllXJ4ZpWZzvzJdSqJamZwCyHe
4SbR2RJ9/SQ+hlwGNVq0/WWtAAGhwloVpM3IymtQ7LSOcZulTBjox7UtmPcJ/dR/NX9BQJikiIJF
UfYeWWGS/rj9jd0G38aMsUs2mCwODqtKUXp7tn7FZlhdBoAO5XLFWlnpuj97+jKMD5iAS47NRGSz
xB2GsDCHgHLj2QFzjkD+C+iw7B2or5K8CFb84/jAUi6w0peWrbXNsQwi5TZWz6uo1rq6Jd4pA1Yj
uGk8GmU4mBNiFGHBfR7qTIx1oS52FoZD+IKgGNedKKmnSX9IczSQa7YYpz8LuMD0E5xmSlAAdpw6
st6Oi5cCLILRVYSP7B1nLn2xX5YFr8MotU+ZESFKR9MOTAxIE/oQNT8xvF4d1eHljX0YAR3yREQv
rCinIHdZSwBMC+7w2jKKImJkA7Wy/KtuqYjVPJiL0EKdXfp4qce0G5miDDDgsDXQoDlujQdKMErk
rnFNoizhr3rcy8KvKvXsAIW3F0OOMqJRFqPvpuxCOppbS3wrp0kFBI34s6xGjohAzmMVGv3gEjS8
sYwUlp5X6vUYXNrP+2KYLBCN7rKbgqCuy1NmjMzB0St/2JDs9IxD5GUERI4ah30FVllnxh2oNkVo
AVPm2ZA02YOvIfT6GcYKiB0FIsOQ3E5mcaaQSTT6PeosCwW3h8SvjClJiCrtk9+iN/tu9FeBc94A
VWKPKk2NUKGN2RlRFexA6o6zO1iiJ0S1etwu8hHkFLq+dOF++2AkyL78luhAAgLF4UrcOJIHZ3+b
sWNmX1yeppy95SlzpchThM3ewJSH074Yi5Fdwzs0RwrjGWx9ILAFwxwdn9UuoLSFcb5ML7F2Ww85
C2sswJoBeKmc/nIR7UCP7Kf1Cspg8dKKwPZjC/Hm0yoTv/EkystQlAB4tF0vHFgBRgZ2SMgNOCja
G36GqzZRprJUWDc/xsbqZOSymvPoLsJQiZ1gKHZi+qUIx1Lf/BiX71eQWDvE56/Avqzkc+RwihE0
H0UsMaxFx21FcSawExSTFIMs11v0AhXLZxcIHOERfP+Or3U45WEm7wJlBBp4A+JgocrelJG4KCWV
70YsZtELdC6uiVEFoSgmgzJB5L9c829lvlJWFp4I/1rcEersMEPP2MDsy48RbJ66Jb2EZatyHsP4
AoDpZhmnL9ucWaMKUa9raPc8lGIrK39DN6iyONkYxVCLF+IBcJGeNcJHxmz/GLsULjbBDWI59QQw
KHS3/7WXP/wstYgsFcxWDElIHlIofZAz840lV8pFQZqqz0mkIe3I4J8wO3iZwM8WWAkim8wfE0lK
+WI19qjBfWQZokAs1uPUrNMMK0mH87oL7kQ47S2xEuUnFuosIt8NvMZ5TtSHcTjND5RLFIuDFHoT
QZ+G8xQMFmmtOAcLbTyg4Jc0RdM86+7rDYZARXsmBMwtUXI+qgFLGBjQ0YmQiRB0DFshPaLTiJOr
wrlf97Jk9dtH70IEkxgTF99FOrCQgfpmO5ECMQ47r2/VxfmZ6c6177ltzv7zdCFznW0anPIK7h0+
FwOKxoiR8Li3/5cQxtNdCXrhcuZAGmfYfJRJwP9TcKj3M6daY2JbwwKbEhXlM4FF5UaYQWQBHBMp
R2mfHh8g6poIM+lkJeD2yfaLap3roQdeM+Hb9gVoNn5RURn7dy+9jukZ3FydTpNJQkMTngI41FxQ
f7ImN7V3A+i5+DJfOVdOXAh2wzRIUdQH+fbHdGPLM72uIx+5w0ZRnIh0x26qVzVKuUiJUGyn8TXF
7z2uqxLdsKOCxqjXhS3eJ7kNff0rmXN3ohiH24tnm4PcsdXKmC5NKa4QXRjcYpRMmzJ6NVyI6i0K
ROwTPyAugJUbU/EKHqRtEzKSgbl58JYzgACcKBrBCT7vtaT+bp5A/ngFcuZhEo4TdY9baWiP4BcR
y5sT9hGuIh1K2XGEu0jHdMY/3Qjc4dNzCcJacyaAkQ1rGji7kh9DMIZanJdByTZZDwNSymtonecN
ybTl66qVVoA4eP5x+rkI94STXpWQdd6iUPwHQsH9k1hLJQ4dKEHTnzoe5Z3N6eCZlZRvKcVbaCp9
6B2Dehc6TKzKW+zkcy+2vPLaWCr/fAXYdmpPMqVAW0qbIydFc+6zcaqpI+OIfaWb+ZmrTp1bqPlh
bnQs6i4Gg/FDldGuvlyFMc6/2mNwGpQOuJUUsaUDZXHPq/lNwC/3tXhdFwiPBySXZic9V7Fz7Wi/
oh5onyGqBV7KYEETyWkCxrmDAAx6dTOlav9IS/E8/DoRwaywoNNY+RToPCKZGv+ZrK6CSti+/skl
C/OCprXzzYNHY6A3WiT3Z7qqvvSU++GL26I0SL5sLaTQfKHs33rh+bxRA9UVai5SxFEv8PUeFU7O
sfRBit8hPuxudVjxgLln7kNvgoS7JfbBD/T3aH6GTJfV+Mv65y/ZkLHyLow4YTEgBt/G1+/M3ktQ
IxIiTSOtKiPbS8IhbuBuEKxeXFgXuHFqYJrnq7EC7GjbL8lbVfBgq0EP9pkVow576jTOPLDsxp+G
whVI+hSwRTVhfHBjC7MLrIYj6kSQ7aiDd4C03esHPxCgV7MFuk6fbSpwTBXVBD5WES0ByGOG94p6
uCa5fcG5ZWnKb1XFkTFlaqgDeuyHc4RWH77o89KfucqkgBO+hPNrHp1KOPrxpzimqnt3xDjCYYwb
DAXEPA/cL/LAQ6B/3nZq4VAOwShz9V+NdgDWvNl0gfmOvheIQ9MzE6ITmR9bGJTROPFbqE6JbKgv
k33NQweddDW6RPwT2yRztDkqcRJYdbBRho9iFMwsfEBY9EEEDZDd5uUcRaHYmHu4+n+hEkrWG4GF
0DStGY5oJG9wx9OEi7cLKcfXpjEC5KYB/nmcmASJpjl+42lrt8pKmyM/mbg0AJAI+SEkdkxz+m/j
M0KUn7ksXasGQfeCdLaGHa+uNeZ7q3Rjw69mYc5yQdDPEF4dYpegpb/mIN8LjVKfrjOFtuz99PcE
1lvP/BF9xmc1/lfncqDkPS5jx38Z3e5hgMB2UoVp/MZs3VKHXj5Iv9j4+I655e+IqOQSoCUve7KX
BTCBcl4gJb8NJJnqindQTwdiTTlI/IZYo5Uba1+9SJaSrdP5OjpGYhPG2nz7xpemmPsGxYxMEP/e
X9dCyvirKk6qRhxJeEVRM2iIvHctG7cM7twyvHtu8FefjLHWRGOawKfSHizphA5z9A9cbLdQvdyl
F/dpUWj7vpRHJMfk7MBUYBpSkeyme5xBqHP/DMnd+IsaH0iJaUtD1znVN//R3C8i55A6dhnVqZ7l
XfE41nVsrD4SwYZAJloSD3PIg7E/WZ8pYYXweUvQiB1l77b9V3xJ9sFzekIlreIuyUphx9b5O8xm
8stDfqUSWjFH530HlWV0iB0YIsCPxnF1/7MySy/YZv5YxnKugscP6gblgNUagdIHUd13Ka9G/2P/
ss11ihulaBKkWCXzOluaptHtk8IhfYmHDlG3WB6EZY1qmm8BaUthTo/ZU8noWPl/wEr0AbLrK7z1
cb4jF5S0STmzuNh+mcChsYLGE8uTgaBComjdWKTl2fjcoNrPoNHlMM2LCaj2+7335OJfct1TGm4G
B330Kqx5NTx2wazUJ6xXqO0WChjhBTYZ/EE+JZc7MxXy+4+fAuG0c+tGWP2/JqahZPEPTKUC10XL
xfMIYW8s+ylAonvVbQuaNWYRsuDpU8m6gN6iRlhu0y21FgCGhZ7IFitmrbynLeW+JwhnwXn5THFR
Wt+6Z7ghV1533hjAXGDYC+VLoF+8QWDr244ByuJZeAdlB5wFFsFfBH8+ktvZU+r0hEYingnIrC75
iSqyK0MF0O0isLMaH9+B4kPn3jrNJE2bD7NIBg84PVGczri+zPoeyDX0SQll6sIVMYu7EaT5Rck5
jVfSWVqDNNFMKZMQk2ZFffNHrPwmdtYGKhZo8Nu+dNBbL7yomc+pIm82DK3UpmhK4K475nSUFCfL
Hp7rV9xp4ttouCOlNH2BlH9bO3BItk0zGwRXSVho3f+PmSGt3PaIFqqRMtX4VWwU9memLPbVlggA
cs0JsqmgEbUFgvfbwji+WgClcU+sE6h6wS/kzF17oZxO9VwMiCNCaSJM78UpRXEUt5WoKi3KfJc0
MtvSXW0UcpRkcUgXqishMOYCW9SLQT+pIK25sAuW/dSgIqZVYuzvJPvFibFa4yJuMhKwpXsARI6U
Kf79juzSU31usONDypMcxD3PDx5j/fpY+BSewri57OEBS8htPqKtC/uL8Irq8qmK4fsbJum21Vh/
NtRLNq73u45GVfLQE+F4fNZLnOKCxDcOKonSTFTEtTK/q3g+qmz9wi5a1TsQxfRVIIuxrVTwqh+a
DNTL9SjntpMAZ6Nfp/usaWWXU4SK6FYUO1M3JtFHlGFKbX2IknJJPqZyzqB3KAEtk6so6aNd8Fk3
/r+fmLCYF4jNZqd2zqn2bOoKw9mi2QijCEMTaNn7FkMNZpadVlFj+LgM6RCyr9ye+PJu+bqrXNgY
m9Vzb9xBYeweLcgLMGnR91rJpxP0MdCh5CkeAq5j1pVexp/Tp0++mXYWnnmSL9HKVnZieeehKn64
eXZalu/IwEvD/6/PPW2L1AganVkwb95ehff/7RJCvbw64HknqrSNQBV+zr8iVY+DF9QK7/VnklAT
u5EQ0PX0zEv0kUYKv7amg5tqrFw0LI1wLi+BMw9UIO8SiqKQOUnFi+QF+mOk/y3XREP7yRFWOqCy
8tjiss/mCaUL73zj3gw69a3n5yQaKwGEOe8g7V+5oQVK/Bn9qyiVYBQR6C9kXC9P/ZL+hDkvr+CL
cIO7IrSOF5ARDIAZJHGdZB5ShzTW0pbH6UYLCJuWr+qTif3V49nfTmPUlJ5ZcG1Zy/I+0yK7SvfM
by+SZdxnavx9u30rA+Xl0crl0gY/5Oy/a4yjQ+Q/W37rSAFtYQzpQlrd5DiZsVoYwRng/pi+Qnny
WlmQ+Ah9wE7+3drThuMi9eJxnR0hE08gt/aZKuFmak4yEM+un5V0gBSQw8+vgypCG9k+ND+OqqTF
LuOiPLqfN+rTyaHF/TAcBkjkinm/gQinq56KMitJzG+zfMOe26Ezj2cPjKpGXODSnGwMKyeDBpHL
6LLgKKgO1WFfsJILWG4UJlhHMu8ilovbyp4NQVZc2HqczlpQ6i4JfhDMpGrxKzTC7lOj4Q1TwQJ8
4EvJCny6LLdglPb+EFl5tRSQYpqEE4Jkk4syyUGlWM2KcyxaEEEmZ5IvSrIz1FJRWpLrQSKQjPx4
BxHrtHPDY1PEZ4DTebJvB0Dsk+eoM7Kc+SEwquLLQ2OptivlpBb7d+amfL0BgLuxiaiTcaRtZBlB
RzRsmq2Yng3HDkkrDLVxcy1fDzuEq61On50FaJDcuESlmKMEnY305pxr0NopveQtc6bY9fluXyy2
00Sz+iWOYo7ma41BDpYWmZrVCxbKijW/Hvw3JaCs62Mv+dCu+5IAcLCNNb809CavDHHAvyXgyaDr
3WVqxFBEsXzcyldNhiwXi15bNcBnHH58PtzfsQDSipycSwWlzkWGweQ4poyK9CBoXZOLGLVJsFKS
zchhxS1xqKb3nBk141RnkaFbhdnMt9RGw2e+JtqcpWi9JiHsyfpsmENQvF6yciSPWY2/VCz9VxBn
Ow8/SZIdLhtdmkKXb9iVdTLHXjHg9bB/01fh7r5nIxJfIn9tGzfpgKgOu3WmGTWBA+spsTaAg57l
fiixQ+5esj7MVgxXX6585HDtKKxjYFe493A8unBEncLLnvTJOEdMK8oPzTtp6+gH3pCilgPyRHfd
V8v2WqO0vpG9U2IgxRUEvnhnItY9rxE+5Fo58TTWwoFDZq5/iXsGIVHgVaPJn8K9Ewp490tabGn9
aQUuLjciC/r+GGqnQnADA3bdRT2ycuWMCYTwgMDDA1COuHeKTegUtJXXKmEpBH0IZXOXysuLPPUt
CjmwG0+VxpOjPtHK9nJ1g5cHR78KLrZLidgSMt0UHM/JuiqbQeRdDtjInNeQfczWSM4jByhEd7vh
cR1JZhvRzZxGGKgXPD/NECkeU8akQyX/E5YILYNjsxBsXrLIooeT8k9xnDZumBJiDuQKxBmUVnLN
EZi2te06UJf28ScMqn6SU8+C140BWSwf8Ui2DZCRC4jogjZ//iRj5aEYLBx7w5ROKToJem5IIEZu
JA/brN3/++NeyQ1nt3fdRYOhHMTbzbcLSzkSySg92eEYoSIG1rK0PEnwWwIBTo6AN4ve4ltvjy27
ZpnnrRsQLzp3TpIR3nf5n2iMhTitJAc0EVaFT5AP5BrB7M3JEn8ML59MXeROt8bwr7IuRBWai6st
KpedYyppX75Zxo6p6sHocf6Wlf8+oJ2zNT6mRGejwPxVPJzNt57BF/6JeNdS7iZ4ZTr4CCfBUO5e
XCyqciOnMUK2zCkFm6zMFDBbb9MwaQXgPaK12KajQLr+c+rpgVYEp41MJ6g3kzHb0tM4EKWBrHSb
9Vq/r4TYzgmSh4NDtCtsyzvfPfkLoKRyUqjVdHv6dK5r4EfW/aImQOsMHd+d9FOmBVfWtG2CkQaE
WyFrJo+v9rv0mIZl4J92Vuy6dmbpIIpXQDShldkOtAaWTDGcln+N4AmiLjNpsWJX5Q5LnUXUEIHh
3d1gxVSeuMxCzxpIQwA6Y30jMwd7yac9iNtOUTvpBGsWW7Sy6L6WH/Y+dBjjqRPrcZ5TQI6uPmSM
m7jzeDdDJCojbXxLCK1QxfuZCpg4uuA7GafXRNywDHFso71fbvGABluoOMypJFsAF3YW9NXb588T
VCav1uHyafoUUkM21zJNwUYpkLdcNjg4tDjlNzQA+GzS/MstxQcUKzJDX3MfOzUHL0zr/iwxFCx4
DiuSTpyGqsNJDvUo4G+/kdBeZu8MAycg6xeBl9OT5YxO0Kn9+5moz26qqjPC9HPFMhlVI0//A557
Rn8xzry9saQoYhtEFrXjp0/PNSZIzg7tJtWFT1H0tcy9oNuCyyRYcljK/3F72GmZNRBd6/QWGis8
Rb6CpNVXEyFKJXzwwvSNrAWMrMIL5vSN3IsE+ihhjExaiL8M+f8xVAT+dTU/ccC8lVAxKmfYNQ2+
6AS/IrlcvSGtMkE6atYatGkpALz+t96660SsR2+KcZFANTN/br2gmPTO2RZEggbTVEM1PsK8IKHz
hJz6blZ+QowqNGj1j8c7G/THEW2AdAYj/0TnwT+R0qs1jeXtqAlXIusfEtokt8HTvhY0KvjLuUyX
OEArFmeOVFacWbwqjlaC835ai8GuddUwHwXkl7Vz46KzgeIEfv2QeYRv59QeeuciO70ngBKdrUcr
t4Itao8KpqLYT5+vPR0rmq41uKHRf2PHYLx7ogoks4kr09rOvOPKMBRUqceje7U5QigXcRIZ63vf
z87zGEHO0g3O+vfvjLnNPjmjeDnWh6MMYeQF8fzWfT2IsCECzaeaHKpsCQRclEDDHsPzqoGZrb0r
cppynqLR1Rs52P3Fi3U1arI1UCm7dllrzuspLzm9DE3F/NHtyS+GgfD3EcEbPKIOyplIe3WYCDBI
RCeiRf+6vQy3fKO1WL+3E9kgxzgsyfYU6Dxrd6ks+QUgffuUKz9dw488+yuGTlSl8G8m4Jx+FlqM
HWR1NXwzMW7TvcjpniCvhJ5ZDnLl2fa+4o5JvPuY4RwqT9eCTaqHzXM77hEJu2ltT+qHMJ1IcNft
6UcJ23AIM2clq2+u5FjrwowTO2W/MxaiibK3ErZIATLyiSA1jR40v7cn50bR2QOerYxpXN1f05k/
d/1+OKPVCRALC7ZBtpLZ6J/C/E3YO8g7vs6EzoWm2faEs71758WxgJzxZZjNV2N1bULk7vKCXDw8
GX7gcvvJQMlQ5WepSD6WBYjmvum4EmPceqG5J5yPgaP6413jjRsFu+AGiZ5l420XV+UFRTx7+LF9
yXyywdoAxm4MYB3NN6x6oDH2Rx0VgllSbMmWB3D8P4CJSgdO5OnJznq1ndKmVDWZC3inqkHGri7d
gQemvmlF77hA41o7cgLzKtaKANWvlJpObVjd97K8vkzolKFKEizPvaPRDl+73aW/gQ4E6VMGTGys
Drdadjgqd69SY/HYc/hDcdMJBrUn0nWkVwMmoQyOi9rKzAzrnnLtyjybtlA3k56z0weI76gE9QzF
oMV9GNoznjNIiI5DQS+x6h7yfVKXv17aVyvwdnCpyco7YyfPbLDqBZBVAd1LedG0Sj0sAzZ6EVhL
qx0oqExCRc5yWVtA+nGeVDKwppvOtWI9627Nt6Sfik2Cfv3y81fZAWhQQ29y65/t+8AOf2lc/IBX
REdq9i9t9SyQgAxDGfTjUAsoVxi85h7yE6Ehdu3zOD+JYIYKSwuvQ1bZRVgvkOtBrhLGilXLBE4h
nrrCVEWdZd3SdY1gr1YhUauZgaL33Yzn0qlz46JJqwF4/ogdeFHi0N8uYI1u9wx8P1ne4gSVQrjZ
GqCpoQnjL3LUcrZbM8SpdlCZUlYed80aMDiH4TnNPeIJaHvPZizWvMnH2zYuWnMBeS+h7CRlPsgq
nCdKZJxFteroZ/DDN7CF7GMKq/6gZfvtVp7RXjGiOqVG2BMrFGFICvYiPbJKfREqI1kDvWXkFz1o
uXXFDbsCuJRiQ6M7/wz1jse4R2/c+upTYxbZkx43EhKN6/X5ap4dZmjyQ6Ua/x1cxtcbedTjyrlH
l5wCIWcwlRxNtHRIQPckpT8JIkno78fI5ozhys1TsfZuTAWFKrxoWPHD3m4iJ5IEFT9mHYttV59h
2KSj7jRgHK6iivRmzUzoReo/iEGqchPGIAJmipBh720cvxpXtXITDu9jrgqoetmjIggXXBG94Jsg
fOogi1V+pW9u5z6qVM6UAscxy26hu25hl75lHULP8NigVzE4ifmaZ/zcyyxrKx0ZLCfhKUEYtSCY
tO5sXmSyzJza70yC/xev5vUtdH68Mro3er2hVHbvDUAbHb1nYgQBZ+YslvaGiAwXG1WlzWNHMNi6
qsTyDetnS7emBQ2JxKg1d1by+RyaO1q2jPDh8r3VfSCAw4T8yyk4KwnYQMKkifKq92UBAGRuiCsZ
ZKBu8N2MwdTHPjucKl3vjvMmWo6rOO1drSkxcAH4tv0jEwBCem0xEENOt3me3xCRwIYwL7I8vxmP
temkYCIFJbCgaf/O+E62FQV65he1ea9Pvmwas6gwrhzl2NkKiCZVqsOaui6nafJuswkvWthUk9ZK
Swm1rGbirMbjDyvLcErDPNn7dEiPlw0zPHG8gtzRyVtCgFz+Bjxti/RZw5yqCfVKVTlB7pcK2M0o
89UG15iB59cgonCqka3QDNSx64pCz7T5LSW9LmVq0nudqN83SRKQfkW001r7uXElmXhziPLTive3
yG4O5E3oqvk5E1G/ytj5ChSGek51dnDLgTM3gB6DBKk2YMG4Sf/5qJRc+8qzfGgBPUgeo4HwHnfO
EyjpxzdhOfwBCDMxHj0iDY71lcpb9h5gPp8SXrj7d9cV/tP4S/D/RIwh5wWoS47GasalC9bq40t5
1D/t6EW3rrbMsf3ZzA8p2LWasr4sDOt3WyinhNrZ8dxjQ+puu10QfeCdTHP/QhBWWmVjdDMLHH7s
0C4SKF6hiUjANi08Xu1aqPL++zFQ8pUT/rb1+FYfb67L9fzM2GshWd/dffiAbNVC+vHoT1C/IhzB
UxdGCXD3Ey+YiBC/wt0mrjXwlelDL/O0vqigA6W8gsNgc7p7DPCdd6Kv6DuwuPNYRGOUjlGk5P6d
77m++klC4FrGKE+lU33f+BHeon8pJCZBLSDYYd05/omYdngqgdovn99YtiV84B1fr43XB0skoicD
6LFqKG6KdRldtrckb39a2DZC4//JDz8VT+e1lYN1nTSe+akUm6kIxzaPgsrH/wLxxrFb5pa/Kw5b
TgQIcVIQRR9kN2r8caCCvFqcmBlKOfEg5ithjPi7kfikZQbnRSuGgK8vKcAdkEgJK8iMZdHBaaOi
vzdatNMSWADJNxETwxvFq8RZnfqr9KNi/vVa+uKTRWcfu7xnvcIsdGrHSP0PpHNM5KY/9TCdsWcu
1B4qctZVgxzDvSBtCVac/IHo7s3+bIaKwqHgGpeMjVlmX8sXz8UP2AoKUymG/yM1W3GOvX3MFhjC
DGEEPsVKYQNFjOZ75fGVL1pLjefHloUBbYkdVPGkFXF1++59O5LqYcdADWFIPfW4UjG07b8QdavY
rx/ZZckjpnI9eE6SfXV0AFlMgvwAlnonYKiNG4eeE+CUS/OjHC3voW5+/EFqHhstYlZ/pukp6CwY
GdPzRVd60XoHcCtinJAMZK7D4Laxs1N2e6UKG5qfUAwoBU4U5f7rPtFfUHevD0m91Tzku7E5JXVg
PSbVMre9cEBzlV3M7ddU1441jMuR8IUdwP5HgsKf+7gsE3DOoRCfqscVrUZQIPe2z5n9pIgbewOm
lPT18VQzscuPrWyMQL1lN/XvKeXTU9dqz3Ul+6F4Mr+yno/eFRjQXldndL0lww/DrKEz7iRy/F8o
QXu0n0awwvSl5/i/yWTxKQF5sMjmkZ9odsbwuLrZUMsFnePvbdI2S+dICMn1qSD5Gx/W+vw6pb+r
D7HZ1mMCNacaZhx0aWZxepVpgIafSnw/akkFO5PVvkeqS2NkTByn8a+Mkxj5+xIP+eodskHHHHdN
5Ah5e4eEE4Xwxg/4qS3vgLnxBOvtSETUQO0pOHTmYnUOnhtxocCSBJfYprra6e3/mOsQ4Db9X8I0
KtvF0h9vSK0dlxZh2UpH0EvxNObqaBPEgY+QNKa6aUJ8/JTmCiZQURlfQlXdbGZY7Eof49KuN8hf
ZTxxxsFFXsV+bZUf3n5o4NA4skNuoWu19JbPGuAjkq+fUzprq2QWhHOEbZVCOjQ9DGokE5TT3h9V
CaNfjSPiaFxJFrgfJYqFP1U//cR+a0XqXeVDlUE87FVP2tzrwTyD71Yya+sdADdz3BJIvlQGwgKZ
FvCCN2h76oQfxEk0paU8Y7t+gKPcz9jH4DuKDpZtwwEP2BOmWivDzMIdpplzQmkRjdfDDxMRjm5A
l+ULgZ5hXwcUrunp8oQQPfOyWFEHJ6LyOAk3qRvWANOYKI2rr9qrzJVYPN3eomKHYv23smQjdNye
/Mp3YC8A/2HWAAO5cgtE4MoEosc/QlwC3pA5ewZq13SaulfnJ60XOid/fMYEZfFKMTRrkkFiudxA
rKxPTQ8JMxuwmePTy9f7vSgPNTcgrOpjPcwDrDhRPPYDl3/W/DAprUdVlESn5EO6tlAELK8kyCJk
syPu2MCeNTQXl/W+u3ioURuc1dPuEF6AtIR3yMpRkwAKso7rDEXe8uw0mZW5D3Foe+0K9yFB+E/q
c78LcC2avgt1yvlTdwJkwWGfbxvbXoxoM5ABGqzcjQd3H/P2/iO1xbIErSrW2sRnQmGuCX/eoO5P
EcrHSCA/KP1+E60AWvmhnYzQkcn0M1nbvLbEIH0C2VYN2nbyXJB/RWm0BDPmZSJgw4xnqfOyXcmp
ku8piCQBbDnesNUSQJldjj8RhTgJFaefSWWKRJSZGZ0tYZmUWPwRM0GLT7e/c6JqzXd188dc5p6b
P6emNMObMqWwKX6OVvdLZpOn01kG2PDnORC5k5+0s3Oeip1F/YBiYzc9GzxJFWkCi0AyOGH5z8EK
b8R32vK5DHpYSujk8hR+c2lDTOOiy/1avDWR5s7mnEKhCn+fwEaNHkLwlCIGSuVgYHeFBgE6eXfV
EmHUEs/diJ34TYqjHs5Shtej7cwvmD4G7+X9eru4lRTaFcVp3HmKb3nAtbZJvxDqIH3mkGgPt7S2
1s2Lm49QlPCm/QBS0n2hOe+tk1Dqj/4AN5UJSMXgla/9NVazrpBTG35JVrKu1OtfE2KzdWY++838
3d2CotzjexHaqUW3fz9dZ8gAGZGU0ieDdaBy/1Qw2euxPmxAnN0Qx4d5xFpL4Of7ZvGiaEyew56K
X6ydmzBpuEPtDvtfj6TCx4fomy9V+75xiOYrVpcD0rmKDJHKoBNrP2HG4+EkgD/UDDoB/X7UVs0c
PZbBINZ7AnKw3MKwl0Rjqdn8QLwnqtgr06ngKANF9jffpR/pHOf4PvBwwDoUPI+DHJ1qvrkHt4A9
eRD3x46jbbiZecDrQU0MmgA/KirKgeSy3lSoan4rUcW+bjzGIRX1Rwqte1PoxMaoV0gIIDddg97z
kfrj/DeSb0P8CbfY8xQTSgCdjkXh1KUWCYAnJeBLKSMm1nklpC4yWip+oTemZiLI+Evsut9108ER
7EmmUqjFfxLdYzv/nV1eNvXRIHIq5NJqk42SWbRrn7QmWozqmnRVnGdnerShlVBPAQvGFa7R6wxb
7TBrcH2IBwDSqAEnulTRbSQL1p/23oyLtcZqkHnfy2zfvu20LG5/dC/krOSlCHEWpLGn28SRF+j7
uwVjLG09K/TYNE02M4m7GR4x787Ce4LFXYaZSPF3w2fetit2o+GgFuzbusPi9q7JI0rtP35GhpJE
XkSXkphAG46+Ln9dwgUilQx5q8AOdUtsGJZOh+vWAGfcVSvph+PBG+gGe5G4ZCOb6bu43vC/vDjG
0A9SfxXvO5AdB6FUmj8hc4eNYdEmsdu0jxEt3iq5fnSI86K32SK2tyQf8hltdSzenu71l/4XzLKI
RIMwKM5LrzQ7lqUXscCzcRCwXjz73qLOkPcvWt3cwFbdCdHFI5QASgbKfvVWEYQl3OQ/mZLoAv+S
v1kOvfJu3bIi8L3JJ3+17HiC303ngqbWDT0JN4ljRgc1SNYkB+FI0rvZyRrRPvRwOMSDLRCFwUuW
kE5gGC0awfObZbgHKl7RokqGIR9GjLyunXwu4yVa1fVm6EQ7jxmgYXCabQh2nQhL4OvrW66pAj+7
vhAl8nqHwQu9HhyJBunvxxISuS5IRVqk0FyP5t8fb3BGBTmmrEQVhSV8LGT9Gheh7izt1caz5eae
ApccmcKCOjK8eD16ciUN8jT+WVomfHTNgftNBKNvC1DAEwdh4ZUpgq7VLkeXw3lXujGUmsoIiUIQ
FGWn3gU4c9AMUf3rNDO2FtKdmgo4XK8BfvlCI9TP1/qwaps9h79UsjTV4SeMDV0Wt5knoJSfDskv
xCn7UvK/+QWL3/4qeI48TTibbBvDHalnz8tggIrboupZGROYVrgyecmSLPIhjXu6Mu2Gn6Ndtrur
mm99XPzBe0I9+Hf8UeCnv0JHmzUddIxs21g70IbW+M0XdaD52YtFOoQLy50dINiYhj5PYU1lNkpn
PzI0BeKEfWOwXf+QI+ph+G8IyFeYDvUyhGWTHC0L1hTiq1jmr1vB5dKWxXc0cZ+9q3uvCiRkTssk
pYfMEFaVYtQBCWMze1pskyTyShgMp4Nt8peUF4WNtcDXZlayl9S47KnP3F+Fn4fF9g5qLPX/8rhq
bUfnJwxvaQ2rt7aysoOupDLQgprAkaewuwbAlTJmEIdIgtxccayaEOSZFa9fM/KrL6UNEegeLNco
ZxY6JobfBlGwMq6tqDAutS6qVDApzl0Y+0F7TVUTZVuEP8ns5ZNTXT7sm4gPKoZrTNaVJnLcI0xN
T7Ie/ZycpV7MSwXIeHQu4ImYi62mSNROy2Ku77HNZUFn3MgU2Kf/5qdMNECw9307Drz+EsHECG49
dvaWID1hKiMko6MQmY49WUXoHtxLuoLtGCKzTJalXk7Re9eVTrIAmWX/5DV21+1qf0bcHAzZ7tdO
9DM+FRBPf/hnC7S3HfyQlQ+wgxpne9GvDCUGG4CoMzwUryXOKrlNbXMfEVzpymvIESfmDCxvdJkl
Hnmt7E5WMJA5xBoL/c0OcIFBxWyvuFJ1M5iQfDQheOOI02yzxT1qInYb5aUjh/hB6uYvcNFykM3z
TtVJ9FhG4m9exavABMxgS/6Yza/LK+mM8KRXEdsq2IC8cQcE4XmgfGz0/qa8M6h2GeFPMW3zQKyG
aCgxCNN3q6ngFNCP0MOorGQLanUjoVpJtmmOd3Y6YC/HeE+rWFJDXFAfKg7023dK0ik1uRyLKxkh
Yg2LD/rzYK5Y5+yYasrHHKM/6ypYWfIw7tpvAGo4GIYtED3QhOam3EqxkOpCRMC6Qe/3FmnJx6ug
89xOvNmImDAi7WyB3Pd7MDPOlQPMP1FbNnWRNp7ywm+PM/MqrA4mbhMNyGZpQlVIIZ2pXCyequf0
dAYHfkENe0pMZpBonL6fhAEPIXiDjgNZ2Aj/GuvbO8WNLXXKQ38U+u/8nr80SlLmTPyc/SLl7chj
rSM6kYsHdUKL4hEyOZSg2UABFRjdPnAQ+xY9O84Lm/ZCKHHvNxayzw0Rf9uiFTEijrwiGgCQ2mpy
n5+pvWTbTKEktEFO/59TAjv28Vb5SpIqje824M2JdfD6EvtmOyD5kRYwuWCkTw+UGU//Eu/t6XbV
ehA7oBaWnNrOzXir9JdgMMkmlmSYyVbUo7/Ce76j8KK3boGfiTY/zSe8lTIQPdUyBQVOcZlbeop3
WViS0BSLRYh38JXFe0nkXdAwhLcfAqXHOsZxmSYEJ+UaNDSDP9cJ7YmadIo7/T4ACeP5MdiyZ6M0
Llm4Kf5XFybZ/fJSUeAFRq3puT8dJLsJvxMU77tVtThaumS7SpOJ5iDsPp2jalDa+7XxLEKe+YOT
SpnlmuzL+E0ypKJYPNLNLgEtLcVoT3izcCv6i93kYe6NIpcfbAvy8ZpsoHc3HmZPjTvutHyhM0cQ
LF7TLi5V2fCtUmi19B3Crh1k9Ttywj74RZnNuridgtZwlcGJPkvJucIUUVaaU9tX1nwguQsGD7Y1
Oeu+jsKdnmFlILMj5HQS7gT1Mk4lTDyXDOkIb/EDN1pnBjyH212dqYK56kQzXERmMTg1lV8ni2B3
rOASLrNNac2MXdsoAUi7C5Mqrqubp9hBekHF18M/fm7yXo/NNpCeNHCH3BhV7nIN6oSNQRGOpjsl
wvvfkKdYkF1l5rUqd4wjVx6FQNp1YzsAWxWJ8nFh9FlbMk4wkQSwb3Nd2WbU+/GfJVaFigO6N/E8
9DHOKDvzNQOHA+glYwLXcVtnV5x7LTZZA/AA54vk+SM/8PtaDs9cvxwA1d22zISXZH9PU1JrdN1w
6X1f9lz9xV8hjBe9UXdiFjeir1SWoFZWhhrLjXONNaV/QwC/9yhylrVDAyJ+zHq2z54Wif9ZHbng
XQ4VL5tNXOGQBxIfZ4nxP2EzH/VMhODHUTZ2dJw4GqkoRtRqfFgztA+beQlUoJE40AC83S8xBzZw
61789vx1Maz112i31CelmK8CTyDn4IdgL3Txso0Qc+tjZOBsGjHaFgb/uo2ONgX6Kdc7f32Gssvp
Vbu10jC2MUP10X620kNVar01d4YaXLzUyQW2avqo853NNMbZ/bvnBnxqoKtjPahbW1FXix3EMqdK
Lj1Sv7jVAmTAykMlgkvFJ3M52/dnWf/r2zlTjVYknQRUq8bGE8kIrax4YlsE8Pp1C2wzIzoX6VKy
nLjV5Lq0Fwn8h0VBYsYPk9lA8Xhu3c5Uz9joCFyH4SeShFVeT1gDk11HieuHu7gO+pudIV8qkKah
AvsghPTm5HUshBkBJcto6GhKTZc0cBLkCcpul/33Mmq631tVeO109HBVkMUM87XyBNLnOM7+GEOL
awj1Ca1tOEMbdtOat8vx33PQMWHcBaczDAQHXUZLJa3pilfw2bgOifzG50vy4nHP68oDlavXp5p8
q9tqwDQilSKFNC5uXV+Y8avV+09xtSbi9TM8Pb1UEiRu5lNW4fU50O/re/lOPSkrYi3mHPcOCBfI
i7Dy9mwKDEfcgzEbKBb8pgKW1vGWhcijdLxtyUZb8xffDe9YpyKqfK/Rq7kdvU2o9qX5qNPk978A
WulTNVWnFIWUS23GAgYzzRjGFPv5OczYoH54v+0v1TSGucktde4qqyhXhNsn93nTZhMkII4ysUIX
b5RiniMLf2wd9vXFMDf543+0QtjELT7jZSOnY8vwMljuBSFoOG3vDOGo9MIChy0tSr6ViEfcK2E3
thQlo7qKL0+aZv1SUBz5BKy8ZPYUHvNJfmzV/AhWWlXjG9JmP4ihqIPvTV9nBpaRIGsJfCCLeDLi
bTU8hrtz6hM8kTVAGGQky0qKkqjX0bhC4j1YpmSCJYt/0z+8MRU5kCBn4GwTWLYBH5WmMa/zMeXQ
qx4WMfT7cDGW2ifK8+X1O+avmo9SyB2nHR4mal31m5MdCS2q5z+wEy4I3WFVpmFIRnG0T4pcE6Sv
SaSTzubdN95QYymmBNCodVR9XdK9pLSwD1xJY89ksPw9rMrjJVAzVjjjhlUf46eYWd4UccatayKo
+vp7TLlQ5ezefkOSLqZYvMposTQBedWvp+yhdFK5cfMaEVJJ/qQ8yKSA+5Pe1WvoDIBWg3ZyzzbN
uuflMlUO6xttVuJ58DnaIhGurh/MEYa4YKezK9ohpzR0oIokQtZyNkoOj6lQ1BzWaLoXJhb/crdx
ch0BsF8DVfk13/Gsi0f8DPVfsJHPThWs/5iREz2TmKCPhKNPp5rNQMfWHXD4e+p5OLCQC7XyURnz
5DTnGztH3Ur7HZI7EZb+xo37TOCet+OofJp+uFyxYB14PeTic102UxYoB76mz38KDnIgXml39XxA
mkXPq2WJ3RabMXFvFeKfufujaGb4QcdWado5gbcwySoMQWC0EbMl0IsWR4EFCwnaVwfGWfTtf3zG
O83Jve1czmJX4F7TY9MEKdYX8G5tcrt9xVDWRyM6zgiC04IGu3YXDbtni3MkxaJ1vkymGIBQOt3X
aBfKbY3dsMKpmmf4mVx2xU83VjTQW/7yDnoarDEG7fYks44bI87pWyla2TxBjUP+dyil9TBjLgLU
VbEn3Zic4L7K3ZS8SzpwBgBJ50oquapKM6x7uhOXso6SIt0GPAlO2pIYUU6qjXdSaqvOe2S9Z3GI
nV++baur/U9hjI1B1vJ9p2svrH4md4k1Y1JpxcGlOSMFf5DWoM7OlIL7XGiZTJ4uUSsshJABBxSc
SZJ8X06Jr2IlfqGOQS9cy+3uyqbms26mNKKxSk5qmMO8tOyjgfogKQC0mE9kC+6wU0MQXpiwY8dD
tcxgkSTBRRtd3sjBCTBd3rFm81XafcIsVUmRczrTNlFi6RVjJ/bXSyaIYUtyO5UsCOw9/vt3Wopq
4lTwaH44KvpvXsmSncy9/Eht6Bj0O1kkkcCg3l1nrOnPxPie19pPPuT+WMNiFJU3G5lB3HRt5ziu
ApsQ04W/j4mzJyd2ZZAoAZRsTJWMsoYHnwESuicsZJmmkk1QCXfHC0brz4oTXvbZftDVwP/RmjAf
eh7UzXQEz3oF13aNMvMl3WTSc5d/4OV6OFXmyQJv/pg8MUuWdDHNzRSnCt97Fw+Rfi5QKs128muQ
3jD05I5ek6CyjEENpWN+T5VUaQ4UZqGdbfnt0liFFh2zfPZ1iYAESlJlaxNKwRrCBjzrApScJj+M
Lg895acWQTWjqDYkxRKw7B9qGluA2AZBUZc84tNzklYvx2MNldvatj3ZfS7S44c3SW086IHNURQo
QBZW2mk/w5mwlqmN6jnFqDHwzePd6syJ7aSprfHlk4SRnzHcAuFSVU1f4wLRnPgSVHS56HZ/0H4D
EoIGPj2HjXRU5o3rY0sh0tJEn/zwL7S7v2WvwOe+mCOWlApTZH3Ky27EbQW8NRsu0qlD38dR3x+g
q6v/02tj/NVf5nAY6KBwABLTA9hJ891CLQ+nb/J9HCInCqTgdChwivi/Xdxu6SbDkUeGkM8QEqby
HTiEYAM9hLeZavGbO+hIaLtTLvS2mVTT8w1ydFmbaqOmKdRTBiss5Xy5Qfv6dVewhzClKZAWmXJE
IGwypMAvCFf94Lwamy+M55OPiRcuxegRRUng8bEp6Hv4dtyiTTeLpHcaEINnikpBLEDacS99qr4m
GWvGWVUftDJ/B2S2uwnFvynXImFN0JgDdJza0r+MrgR/OtsjVijyBkrDUkmxzyOLdr8uGoKNap5D
B6yENYcD1J1KJGEbdpw1iwL5N4Z5VAV9Pi0mLhX70b44QJA9MOd1Sxq1mSvzZYznUHrVkxjA2BjC
EesTOxEwJYbT7mtQvYXXrgS5SQGvhzuxS2Jn5rIbxRFzx2ZapagKVlPPt9Hcwejc890/0uRU05v/
7OpVhwhE0WaVbv4AcaGKmUN2CmOVDgUeQy0+3EdHFsYJ1FSFHhOj9ibdFLkv7IL8qpyN4o5vfxuh
HjaGqAuCjlwfY1SDJDugZK7RSas5s/k6rhzMzriJObbWEXarivnQwbfpgBMH0domN7NOrCVhiIJD
surmPNYdsoGWAO51YOYp44Gi5/rwRc40+dJnQWZSfWiLZaHwsHiYZIz2KxpgA1iBCSdDcjYVxU/5
uh0rXLXD5kr5QK5JL30v/8JE5wPinHKX+MI1ccUBXrk8s02Ht9rYyFVLInM1+riz3CAoneBEBa9J
BTzj9/ODzbhpcC6O1dSViWyjeZuFe34dC/5xaI64nPvYgU5+/iTb3oI1Xj4CgGxdwRkyTMICeLgZ
ksvmpImcdQQm4vOOWSGDRExR83AO46oACd9uinTC8KINGsu9S2UGLWmHkdQ3DQl5Eh58Tz1Xo5N9
GOVAHDefa+ULYaV88oE4jaImTkP8cTKZVJTgpMJkvGRsz9atnELa0gVmpDEtCe5OTVh9O2dnfADL
xiShsPns3QLBdApCgym4H8f2b7dxZB1y0glEYZows+h1c5LXP1j3TOfFndvf83PU1gBlSAZwHWvU
f8oOHA0lNR/DvnbXGcBxEDZqUSrfq2mILbJn/YU+un6jE986u/HJut0eQYH42crhpqkFTDzkIWgX
Hv0VpY3cxfmXFMb28Xw8A+qrcitvvuhEM1KAyQNLpH94SwOL8IP3d3KE2MKDuBDXc4nvVPfkLoEe
VfHwNEk9q7uAcrwBCShQLT+7JHvEtRUF9AM6QnJpOvQMFJ005/widQwT5CDK4wiRP4r2Q845wpuQ
xlHMKdjHiJtSVqIQFcslRu01+1TKS3rvjC7jYLQNR7FcTiFvMJjHElh5lgoEFXc+QiJQ0ISIrIg5
CQGurXe2ZE4j/W0z8mW8QSyxOZAvJctt7KUpkT7LoAXkvf9XMO/bl137aj6W4SA6Uv6IUX5KFkcC
9tAKYISHuxhmAJfUsNRrIXSW55wFIFnOjXH2mdpGGDOK8tv4Az2MWCxjo0SjLRlvHTYxPo5EL54B
RlHLNbJ737ZdOnLCQj1VNywLWOZXWnLygKGTKWEcpISdRRViDhNuJBu1/l1gBFAMH8nTzhGTBGbr
JuGZziFZc2SErkdHdOSd9aET071bo2Ji/5xrta0QYCXdA/92dJxqtxttdY1aKC/Wbiowu0B5zmS5
IMQawoH4z16hGLBOXtiBgvwf+1fzzwlWlqL5o1s/pF7OISE5+96zGwzFmUY5bHMY0aGmqVeZ4IT2
JHOooTxj3qG0q3b7kw5KLhn6Zo5erGWMLAD/7q8m6wnqL4MHV80yncsxB36UGIYemnd21DsVpa2H
DinTYLtTHZUp0l4LmwZvIOqx1Ca9dfARzkLGN1BRXXq4ZuOiLxdyqIWjXnUdxbY/9BUotN7LhHLp
1nclHxjMvAyq+RS5+8s89Lyr9fKoSW+qYxxApbx1QfpOhBe/jrHsJ2vpuHrlZfgQA6QOxS6ZH00o
zWjL5Ckw4EfS+uL1uFGZgZlwivRfgP38+RZ4so2OihM8/ADU3HR7YbHT18uSZzHHasecVNxOBtE4
5FTzHSoh0y+wdvQ9lIWdnDvDbIHSQqgjeyLxF0Rv3HQ+Nxt2TgnLldj16oGFmpqJ41/kmpoF7drk
cXSyW88Wbip2B8bIl7jPHU1z9sPvbHikP1tBCxc82zkcR3JZteC4/pUkrIMtZEZ/G5FF82DwAvFN
Bz/usvhLS3O9fFk+4/Dt6BydYDRFYOfIfPEHCePWqp5m3EbLVifIslFwlgNFlPwcuCDt3chLfYE8
BPdXgArLHeYo5Mo+pvXj/2D+HCmTz6rjjR3Lxx1Q2M+mS69h5SNjmiWzNBCPCaLziVKs1zdW7kVB
mU10UF6zC4D29p3YCp4hfGI+5+OG8E/PUirB7NBh7Q5BCSiZVrBKTbJevWHgxox+1512FHA/3VL7
E8wJDSTv6jmRvKZeNRWehIMETTVZQU2MkvTAOAQMYLr9AM8NTaeZkGOIR++f00il3XkkPG7eyseu
S3LAI4QPvOIbaGLfxguz1V4XsBX4Zg66WFDVZD7ycAkTlm2rX/PKqcoS535TDZ2kfCfY57BFi0Fv
aC4+WKkdw0QZ0NktO7uHkw+WXx8IsjqKqvctywUQ+5JldH9GSkWALxoqGqBlVCBc14qLwEqApdDk
2t4QfaicWKhd1j0fvTSSLcuxuobihRNh3cZH9zCndxIAiigE+b55w2/e1Usfyus7WrUpQLMdF+QL
eaF5wL/nJ1zolAuzd27fxGkanuDkZcMRrCXsxGjTotDX/3pUnHczN0XWW7VVtOK/MWPmBHt/mjGO
zJQM7G0Dh0mkdpywynpL5JbxglyNUlbhVU3lHxJQHhN0qHTdyHGaIQi+2Lq7r3NvqDVmEm4ZqFWm
FKrEghA9HkTsWJKqtLur6ibg/gMNqWjTFcPzIjPwkJ13BACt0OstD9+dhANb2wtXGv1cEQQU4O9w
orDDT/wpDTa04fy5Q8NsAQX4H+72LcXVcSjaWI973n6Rum/XKhKpuuD11wyE2HzFCBXe3tVZOO6Q
ZgooEEQE4GExxk8XOr0NKjoUTfki1zLTxZhVhoPukyxplQtSHbPfVwb4xIN1SmWzIDJrnc5OFid8
aWHsZDuNXOk/Md29Um1vBSFbIAhe5ZCmD1n/EEBGrkmwnnLmF5ndiCzHoRAIYvdLFbkOlGgvgPjy
APDnSbbOn7AaosYx+LeNFBreOanXZOuF8Y5YEmR9WCfYy88rWn0Sr4LUoO/OrdhmqN8exi6NmFo+
c9f1CR4roUYvN5gK4UvxB4dzN7KV1+bpapVwSQHI1GFSrhhh4sKi6OuZLnPE3uVjeyS7+KGqC5wG
sic+HupJV0IM01hMXpGWyfaBPJEJmigDsTCGNLSYR52dftPIVc7frN+rK7S85TdGDaTnvzzwxqdm
L7nsl67xCakpp31/OIZfCTpZDY/am1fjEbDjzHX43qDuTWx2C9AuxcRR9vlyEcUyxFBAzfQwFCtC
wWmfsguGdHSmu275axDbz+C7hdtaVuKfWYHkd6hIp1BSsvcDZvuZYs2uEO0adKxVF2KgGtJmcG4t
9WArDy3Q20s2H4pj+UsvW8dwsewboj6W6viik7UoGmXIUNVarO6bhrRjs6rWeeZ9r4jnk4KvOOQG
S2bYspcmLhR3GSrDYY4WAV1odcCnZ1gDrDy8g3+dsJyomP5IAr0V0Dv1XkPSbgYRD0uwEo7+Bwcs
pCnzgsFzuemIq7Fd2wvFt1H2YU7i9IKBn0SI7XjszSzxZCi7mwxo3Yp0rUreH7pi5uJ8P5GYNr1s
uD0erqDceSZacZD5vzE2dPzQQ01cSCaW8hdNSbYcGB2hMMW70Id9sqfgnXFL6eRLjDi65Xd+mcJo
fRmQWgTCrrbh+fw05e1wbdahYrO5c4JSMgCMDgHQ4iOHkMPV2Z2C0e1N2oiAHuOmbV97YJKmdi9X
8Rl8JxAboc9ICXy1BlCi60ORGdztvmdcxBb5jMYxAojIrXApJAw4qIRnR9E2Ymx8xbQwIj4b2NpV
27+Vrsw1ikm+W55JAeuOLMbHki/04xL2Cpf+kE7ToWvhEC5EfSM4kG6PHUD3nnGVgFs90T7v2Mkl
UGWtWANz/66yk9+pwPxK7er9WEM1e7ZgTZikKIL9LDGFFh7WnqhBkdLPzbB3vMcltl13x3SIX/Mc
BOBUkV8HXqCVy5Dov9yln0XxVpaAngzXfn6zaliWfMKdWzBeTsJO7aooZ8iy9EMysD/6CI58XnJs
KZvwGakvwBTXIJ68LYQHt3CR0YTp2YE0bqgnd6DzDCvshpDlfOUf/iMmtdFJKFFQpfoWF/M7LNsO
JM6ULwwyDbYko1QY1ERwmz8TJAK62VbQeFZf2s6/PVkis+YirhUwbUp6zR3HRmkGAYdmjwVRhtEq
wLMUYim/eFAR0wPeZbTlKSzzwkCNJ7q2R8tvCZiqUB1AnI1UMz/miAQ473kYiDkSZH5tTuMbjIRE
WvhKaLSgxOD7nBdnntbbbarJH57rxEMSbbJup0wxOCFiD4ZW3d7kP4JOwjLJIOlIPD8+fPMk29qc
4D4l1cGJiF8R1+WjZqAuHTnVhMJVZxs9Tc2FVLfx4Sf4oMwtqSUniJw70nfw178VzdC6DDXbdsaQ
PlZpezilgxY3vNtG6MYuU7e+R3E2TDYYJKdDW9w3q815CJHh4sUVKhxERLOXzexrAV7z/t5nbe7R
IMYH9r91JgggzNV6/0LMU5WbYOCVLuUVS+wVOU/dX3H0tYSLpflP/0zwqrpQLUarZ5XFlR241PWM
F4kk9JNLlKnSLyp6kWOaWAqPHHFBhhADqvTwK5NARcKe2RUrcaIoxcogKibAAAyuHEm7SSpUzL/R
llVrbJyLBGMSTCW/bOhTj2T92Cx151H+z+8cSNV13rO7UcPDF7jpDEbmRp+DK9fv64TruG3puZn0
nPO4z7t2avmVdMCmydBhQi0pjp1JLeVrJfK6fSv+FOEPrMTuXK1jP5HDzRNL97mCic0gzyiQdYqD
ku/c4hmJTu1qi6BdMSXbxMcAC+GXDbzlHp0QVdNtUSciOgm14nu3NLA0qb13+Y9POcAjHKAE6bIJ
PwhViZRgDbVEXUmRENkMdcmUnG3CXWaTD7Uva8Yp+UP4m1Yvszr9IMhU2mAnlgOqsWMD3vqhsxPl
qCFD3l4R3bkfY2RbEXmtOdqZEU4WDC4a7o2FVhAjyCO8VT+k2A/bzLjaGexmMuEETbdgi97lsAhs
3rAJOMfKTOs/Th0F6EhGgEO2H4qbY+qmWYlWTCcYPadDTnh8N/ON2WzQs2Q2tEAXjYp9ONASXf0v
aC+F8pSQVN+B5N+YhLwwJiVdw3dgLcypojpAYWXArMwL2E4vj1GnHYxDsEqEcTi4oue6F8HeEgzr
+9rFARjuHXDVkHycNMZq90XetAwcv4ZRgSYiP/j7a9aXX6ifiR8qwPxGUVVChmK5CuRe77BeKMYx
/0wL6QwduEV//Hn0pq7dkqbSqki5QfozvCbHvtnpC/nlWbUVfujZOdGBpBJzGmnIG+W+MZkPLWZO
KSdQGVJwA2uvuWyjwR8kTnNBFArofCZcVq+DPURhCLlUpH6X8O7SSE2Ssxh18nCiKk+3D0Fqfjp+
NF7JGfUO8b3Ny+/AZUGjEpEDTRt5d1waeKeFjys2jTvvoGuq7CZRRjhnuxKBD8EmJjoNq4bNDrZ6
yRHvyYtrqXsygibar4bckRxSEsRSAUaM1eI6EO4XC3pCPrfxHo4EX0XHw/IWzdt9iZbBNF1EtYfi
i0CtcposGdh5P4vCCkCeXmKEfdNYTb/y5645ZEqhn5lu8pxFpH0OFQe2cm5Lk6JqKM00Pc/TUrla
6sxdXOcfv+XRYgmg8eRUJSgfhEAj7VyIVMoWoXJ6bqTW8DMLBCEYKqV05joylAj1113jORM6Nnsz
ji7/oX1ojhN6RfnPvcnS3xZqAQ3iCqKYNt0RFyZzXY/lMRVL0vBlq/NP8qqu14Nksbd4kbI+N1+k
7AxHWGroO0mL3Okr+gg/h6RSoteTb/wJAblQVCd/uwwn7R+h3pS5N0lii0fBrMDGUrW/Es+LSUk0
Nca9PtmRSzcrinojGOJLbJGIjFDaUO02DUxeMZ3jAFcKHHbZIuvAqoBYBU7z/MPohjG2vvpcJ0xL
N077N7o9glnKZuh/Cr9mT5+PN5+oJScW9g5i6qmuqk27QyBwCwLWYe8RYyWIJEujT9zuOCm5AoF5
+GRfK5VO6/+a+Kv2qvp5bXDYwSIILlhLDZrQXlLu8DZL92cxHrRUHni1RnK/SFl57G335tz1F0zm
7MM83fvvnkCKOEvUFjsdwNe71LwwDFGC2KBx+eDlJgC5zaVGNrCqe/j4Oj8+c/jrpeRg8KA88JUh
xegjT/IRLcXxi8BN70m7UJCgc18C7Ts9zjj7rpuf8cQpfoB0z2V1MdE+na4Q1BG1UWatO7z9azv1
BCAK8JW3ORc4uY0aw2iLDbEdlxPLLvOd57Juidrtua5T5cXxNub63asvIbnny0c7BwASwX2pPE6p
ieeVd0UeFHepyP7Ebhw9brtNF8W3CryV7Opl+YfUMZT2J5Peq0KoWQYoRFAVDF0uEBoxdge5uD6W
nnLUc4QjLLLKqEeD7GAplTsKaTeWgkR45Jl0pgvZFl41iMmogKtyK6JFYrKSH4JlcJu29Tua0Xyv
O9tddjP685iA3Ut0QElLduPaLRKm0c1+5uly0k7ZtAIen5ZlP664iZ3C0OA8e/Twv2qGY0uiDpzV
JUZkjf1FOayh0/crvMF6i1J10DsObw9ldWpFESz1UQcGzlPgaGccAHzI1t/BRXaCVzPHHE6rwyRE
pBpwHKAMBs0KZoXmEFWLDJYtYSZgRGMdsRriU6/0K+ht5oeXHO/InBRzjesizqeudnmdpU8pYyxE
uj/3B4rBU1aLvOoVFbnMdjRnihE3CtZRFlE4JMPa1t6kCvAUZQrpbexSpCgZ8Yplbxc8cY/0I4Ir
eO30ONNDHe6gBsr3hdRLk/6EHia2WD5/0xX2bGpMZle6BRbedDmKcNeAg7zQYIF58OJhiLmjgVIP
L3FQSKTJc/l7qOPa4hSs2kaXs9EpTmutEgfBhBe3sHrk+y98PKo5sVcEuCoxTyxSJ3i0xEwI58xX
eUGVSp1Ty+e0K2VviVWjBX7yjWRozBsnLi3NY3+PSj61D50nUmw3Kfyz6KrLJeUX6n4je76Uspo/
adtFQs6s1S4DGwRG8q/VPM9DRfaBSh5gk4RQS3Q0dKmwEJJBk8rED/nukY1fnyQBgODbClib3ouK
jVczaHp+vY2NqTYlE+u45vaJUVhsDg4ex6+U6bTaD391+khdu6PFev8dw/+tD7AQBcQnwM0ZFUSh
u5fE5wlwRxzFWvJ0d3brXTat0un9u9iju2WpKSWFYCRFP4qqVXzWxTT9k6nuN/slzWydrZN3ects
4icaVzXy/HRCozYBYGLNUI0I9q2WXVqObCNm75ZGn/W18pEvwQiDpwHD/AEZwHY+udpRpZYLzGay
qrhuMAVEjazzQwPXDevHZz1fwzlBukcYg8N9AjFbur7RK44QGIyGhdNCf3Dc8lywq0qn+Z7M69E/
WuSS9jmGOsHSOgOz8gU7TgMHYLbfYraCaHSPMevlW6kiom4BBW4WTONme6Tf0lAxI7vC+cJUg3DH
sSwbRQDtw4Lzpm3rv1LV9dFx1nTAhsQaR9VMyYwbFE6fR+CD5KSHGRLTsRnnAw8/LpF6cWjo4ESZ
3sZY4557P/t4fHq04b0jhSD0QrOYwjn0D6Kri5hq54Tqq+xSjEJK4+/TY5caZTC+HGGR45DxMQHw
BK98QdA9jhLypvZge7sfHLMKk6BfLsfzLA2+UaJ9HygBUqoVSzLH7a/14bqjSjM4WnR7keLNa7lk
9NTGWOUslGW0hxAQgJDcsiQZZozT9DZTe/MIvKoe+7S9o8SE8RqgKmh1s7KO56IE4xpeix5a2HV4
STMXuwz2vU1qV15MgVvZPh0xMEudEDIt3oJjKHgXh9xb1zJHPfm0JBfitFNVm6TlURIXtKTPqTaJ
OK6T58lRDU9vzVHoxtW8d0ftBbaEDAAnJxZ/LvFrWStCzS/raZ9gGGWJTQ0BE/m9QlhQFu2ZqE2H
nRdc5A/e4RbxoY60sIfsa2d1+xjjP1/ir/912uOBXGvPnke6hIpGDGdYiQn4unuUo45UBe9QUjEY
4ueE0TPbJ7IoPRHT9NIL+KjKYPHm3LmfvU3bpPRRk+pXXR8OtTNn1qClqvoxTJTptWN6e/DK8ReQ
HmOh9xteIAYiLHniHMW34HofrdPdt7LJWOXGK3gxbJFmze1Ijy6/It9AvOMIL3uoAV0i2Gwv1e0Q
RknsqD4zpD/LIn0JRxdzMI4eCVOJLd7Ge1ejhIxZir6wnVc4ns5QMITKEcxAgwOKmEkIfrhApr+P
qFZM16LPmixPu5XC5yYrJ39ziXVZrRk/PP6Oq1v6KqYqOvnFw5C19hIAilTS5O9eB1nFwIVZiwPZ
VBs2PGpcFYtkRp8UlkMwoCLESlNwg1qCWvjsxkxBNCUEL5ROomo+NT6K/sdX8gQM6YwF1njrA3Ru
aKPHZ2Zxu2dtUJbvNXizRho6XrgnPSm+nWUCHnLXXssU451kaUxO/EbT2+83tfIm2UOy54QnyOlC
ArWUyMvxjwAI9MoRSC5Rpbx2+GjKVdSULA6pDY0ez/mjHusE2aVDHTpxmmCRuwYXaGxEJVYWYYtV
z222tiPf9e1fFqxP1YGXI2sVuCv49uQ1/h1dHU672SGTjpMCARHRLb39mnKvT2orBDN0FFUQuv+b
PQbxWFRqIHlMzz9IsKZBZjATAl2QRKo3FPX4o5Uz3mGoOorMMY4RwdSt6vCjJovfQ0OUhQ8WfK0g
f2lJNJw87rMwpahYFkNuOkRi9ubklBts+89aBoh3A04yEWgbutdImVOX8iMnhte5kF089VgDPoHx
DDWkkN7NVy7astlL6hWCPktTAjL/xuTRKkc7Ld7FdjoB0ib/rUjz5ZS/7V1pUmh/Y0LO6Hlz/Ifi
8WU8NFkOnx/GPmuRKaHbBmERnNIm3x3qj4lO2Idp0isjTuHEDPUN2QV4u62hhMNNErEowCIiI7Lx
vpzW4QK8IqxebaRa/KHUFyEcV2uqTCN28ttVYMdb2LZQLk9dklHVhnlc/UYaGUL3eXoFKramdzpQ
gSnK2NptVNN++YRvJc9iTLSM4ONdvmSQ4IPsnItYcGAqI0b3qL/v9SAXj7uSHiGM+q0wRlcXzCY0
KPowq3+nIJi1GUyNozI6AtzkiP1WulbSXrTm5608mlJGHeFWueiDEQAHa+MLNYfG9OaY2pAoWM6Z
LYLge3UIn1G72ET7JuX0Noz0MnVZKs7cCWts0AZcmeE314G5XtLAjzGdyxvSJE3Nz/qsGdLbVmZy
M9SZkEI8HM4JzlLom+xLSnQO5OaQLpT70KAQ6UZedbHpX6MdWmfbbz/zg5AOjGBSbRu2mvtuRHb5
NGPzFoe3nYwbjiNLLYWA9W6RGhhHl6agAHyAInKRz9uaytGQGLSt4vLHvvErg+lqHc2rC5kIPvs0
FWmD1SU0OsPxF65ptxAB46Qu9hmah3dEX1f1Ia2GAEM1MCeRrrrp2aryV2FnF6DyjgVvUiNC/B8Q
+iHsb9FK49h7PBdOr+i0s2xRk5iU9oSsN5aB/tH5eiHpx/V283FEMH8ypyUrJGR7HkYFLWaaUX7d
SAx9Q8QuZLrxSxrb2gCqVhjXtsWBW1My5FYkzzag64hOrKkdE6mutVcF+U6MnvssBVPefBaC9oX9
o2XiHlAezgjoSX/lFYJSbM3MvNLKcVzAl4ZvflgAVWtmDFhvsjim7ByHUZfVdRs01a9QCYukYs+9
AoRGmz9P9H3hOIq/9I3WpNPPziTB4mQgsvtHo9cmPXBweMidGNFuRJMmJBtbsQbaYMjwJkz2z19E
WLtsvZob5qGJeEO+IajH4/FRrHymgRqGe2eJsRtteuLbLloahpJAOrVvet9W8LHyAYC5G9fYj9It
sxjLSN/Av7ExHDJDJjkrLYBCCzTDjm+VwTwHADkd38vPJ7go+gtdgxcpzeKJWMIQ+k0xEgqjlx+e
NFjUTlxQBuPJ7TpsdYUoHOz4jkJ280eiJkJVX5/Tb8CdhXM+3eklp6HrtQylxXfNYXGPv1jI1pAd
pz7uCMuS6bZ1E4FVJrUDvnurxaaCyLO5six7j0teHDOYZ+hYeHRMWiIGK1U2AkljS52M68t2JCDU
TvL+G/cts6nPqkIOhjY53h9c42XXNBSPKz8mPHEuLfg2DoxTTQtmlW40aGStUoBoRggKwQ9PABHr
6gBEG1ONprtWg7Dzc+J9teH1QOIJfntwQ+FT1+4smaKKsC9qElGttDkZvtYvbDEj73fW9lDm3yIV
7rgKYSBZfLPi8eDnhEzDve8lNYSmhYa3o23sdT8UGSZS8Jh3o01OVa3YJgONfVRjSm0o4TvSBhS9
N1PZDaKCKM9YXS1zeBewak6M5aJKWg8uBNROrSIJ7Hk8K+YyoP59O7aZysuHGY2u2f/JmficHnTF
Dzz1XCM3lID337cnM9oFUiF6JHq9K+9yFdfB1VrlSg4PLP5XnUDYOzGxjQj/inq+Ue0Wnq05HVEX
VvKGfbtueFrubxtEHyTX60ciJDvlxDbWzDAhm2F9K5hS6tW2dnehqIjbpFpeD6/r26DetkOmHSeb
8gKAtCB8g4M8hGwZ4CHz4WyUTi6BKtg82Y0p5bAIAUPHx9bHs0cXT7RApgRPCOOzJSsBrVvgmPFh
/9MJYDMpExyV0oSTilEyT+9QyFS/jWRQdFFepSoTw6sQwAdDuc4i8Dsl6M6RTBA5faEk4rG/9RpI
ESzwaXfXL/9ePU/APFSGWHAdU4U3PjedBDJgzxstpdmQzbn+duW6JustmjLaET/QjA5X2A2QVpGm
Jjn2C1qlZZ1AaG9tDJTp+s47WKhDEnS4TiHdzKZ/mSaU6PDmMJzccmSGPMfxbmZkK0rUQ19sN/if
KMb52WE23sspmGqeUtaEdxfnbiCnra+bP8su4brdmPX4JQfXjBKCY3MlMMp7TLBfQ48pljESVJiz
8TzwL5nWzsXobe9IuKxxyBULdARzqMdC8oixCa5KpaGbCBaXXNpnaOer99fktBI831h5WU9vUJdN
nDfEVvoPOxEcZt7B+SCw5y2vpyvtW6rcOCyAdYCAm0wyr6HgfS1daTzkI6HGjbq03sdna3SESsiu
ePyK6q1R27Sn9W8N08tLLliFAYMir7GmMoX1Kbbb4EEvgIT3aVgnMLlBk9g3aFuEs1axbkgEdK9x
91Xd+MLuWBBPiXM+4IsZvKR6re+tdfeDaBqhHZ2huWgjJgCgW9XuBbuyx4Fcdu0b5RyEMan32Hkz
UQz8LFrTYqIGLjzz3qtihtqEjx6a6O76kpYdYsUjhSO/FlEY1le82GMNmn8Qe2uHUkrIkl8clXWx
yTgNWc2FisdQQ4nor7KvvLC2M3PKLphy6iE1LHAmsiAOO+Blu6MfTqZCgHDQf+kwoErU/dUXlz95
aSaTMdlicANM67AvkPJf86C+mGHhX1CH8ReO4m7fmz+H2ECXaTR/G2ZVTA663c2BS2SYSzIfz5iW
svnsM2u8gx1M7LH5Z1SaJ6tIUcGX5XMWKmiRyzKTJRLXw9oXaFdSFnIQ6uzegjKk3zuBr8kXlJfa
xKfIB0V3zHHopi2V1W+zKGzFdsawv6gFMX/DqqqfV2swPPPpA2yOdPQ88Z7uhliUA4KuHsEyvWsL
3hp2a8DDnnPoyk5wcI3YjfK4tAE3y2l8HZNtYV00EOTvrY52n8rYUnu3KyjD85JxojeEGrHMbyEe
iump8mDGhpPuaRHYHKFuRLBPw6xTvf53JdAkr+mL2dgMmKo+dNJSE4+3xkg6z08ImXtWQiWkwty4
36tyk25Y1FPXRHvachuDW2N+PHMlD14i2IUGdcgmCa32blEYOk/kdBtMRN/TSb47ft37esIcmpK7
GXIBgxaExv9D1YE0/gytfqNZ3r7GqV+GsiqW07+8A7YQ+ZU+twmO/0oIXZejNhvkqDqBLUoNJl9b
nX1VmttvrM+Aozv2B/v8iV/wIdxi1W0cMEPr+cOEiozgPqonu8PBPR9A8gtlIVkewlJFRfy1zo3q
sKQfv/bdE7TX+e5qXss8AYgWEb4pBrrH8xVB1VtIlEdoYRD8HATMH6i56xUqjwGudyQR7kVWZRYU
watSjGcJaqtdkDz5Y+xUuP15lnyn87Or9Lpc2MpPxtckudOqM7JfMtkmG9dXmAdPED8GOaho9UyI
u29seWVWA5pAe8rLnIKowQxnGRFPNT2TBgBSv0tD3fkcDHSaOAbK74Ezt8jaIxGMe1iWeG06BAad
+DpsDxWO844W5oJ6BEtqiA38nVBXlW3s0Q96HxMIGKZTI5DrM0CMXr8JRkL6Gv1eTUELNvLsvjF/
piLMwLr07e2LHwa5E/Uj0S3l2wAxzRoHoI42X7CDEguRflEqdLzjGgJzW0OLh7UUOhXVTNsr8SBJ
G7SlLiHoT6rI9NwaIvjKJhCzq9mgM6S8njzNGSr8vfnMX6Qc3c02qFz/Gphc2oRkpezeT0EnLvay
c9HPKUARQApv78shOi8cN48/r7IFEMKIXQccvRCwVHTiK3oMhbQYm6BnTi1akzEOvE6xaJvRtAZu
jNVDbar4GBduGbab49Zg8fCYKotTilkihkEetzu0py5vs3kiLNcAr+tKaFDJZf157uenIQx98dfW
2cCEYmSdsws7CETVaJf1wAxwzduG/4Sa1zoNCw48JossY8A6+ci/eqbs1nmrmP1qn8xsBsBNbfnb
1pdXSFO+RTdXD0vr0yQSsjo8tVtwcquUE+onHkQPqa14pwrW2cAwhWaSjWRTYekGdhyQUlYSnQM0
VV9LgmLdeTH1doiauE5I4W82/3YPLc364D0QR1wLIcTCwrLxAS2qFzAvjcbvktKqga8+fZpd0SvJ
79BWR7WIt14ZfB9VBKlpIcorIjzNPbTPd5TavlKVCYn20sR3WV/DgAK6dzRDnIY8nhP2xZUf5uWS
bob3zn/UiUGhPLJD5TJjlKSgCNeuzPEk9WK+q8Ol3H7hpsbZmwxV3U8Ifk2480w+gGT/LdNy+AnR
zg4lRpD75sY3mFYi8QFAtJFdFZqxb8csDfceTfVlvHBHqOZ65dY/bt0pk7PNheXUUm2CdauDvT1P
Zmf1TEsuRrKRYzLBaS9AVyHAqlkKDR9nEzLrVACnpSGPbwpKudOiRWfd7D+Zt81/Hz+vdYrgIbCh
zbIEWi8HFIYgF31BWsh4+fsozfINIQJrNa3y31GqyflYehuqd0YY+qsb7BsYQ81MxGdZadD42Bah
DBNp9tji2ZEtyNg4czd8G2AWidCPdv0JhCwksX9D86AkzVfImMOrdeiTfSSytgl5D0Hr3SCVBS9+
UkEcqX3dkdigASw+EjAMk5OFTLrtW9Uz/zOWG4g7Q9e9WYC5hl3JaDaYnPiKDvDxw6cbCj0esiX+
fJUnvflf2MFZM+Owax8FzuXKEZl0Sx3GtxcBbifJ5HnKo1FgJm8euYzq1W9WeVKPgTn0/NID3Ppx
TwWchxPVzG1YL0PJZsd7UMiU0AgcYFAN0BfDaIrG9HLQ4KM06Ngw44MbIi/hsRQQayeO0xeHJov0
9wBPFW2lVhcDtrMCJs4jMI9JBQahnT01+hwV1rR44a3tGmZnUGUL8FfqXWCBIAeQLAoFCq8hllS7
iWY0MNWoWo1wW1S8Ow5jpCZZoWUJ0RfSO2mm9aHIvv19M4eZEVS6i1S1zYGbps8ERh+WkLM0A1Pt
lmJn42+/fU+R6fdO7rDo5LBske7vME1mzgH34V+P3tySf/7S4yzvlHnFF4shNVRnOtrveDl6niNX
vNC8ydpt6jFoJywpm//r2aB0QoH7RTIgPTAn/lsR3GO75/rXcU7lV0ZjuipnoTsiiXlRP4Z52Kej
i4JCuotIt81rWSMxn1F9J3ptClEuyz3cY6I4xwVEkF8g7SZWwtrKEYLG60VgkB2KlrctokRwHNul
v4lOCneQDfBMO18yNk16cW7bItYxovLRVADC6yraBgRCsgYVmgMnTJEL346AYVxWjuHqgKSFJ0mo
uXkQP/cPxiDbmGzYYqsP/ZbtRStGg7m29F9hq6g2ZVo68xjpcWTni0jZI5No0cGlRPDzG0h1WRj+
7SZxLe9EsXj/6AMUOz/AAFX1sM0M6YO9m9pliFltBha0K53H3jkUorvRYY9GZW5LC9H743qd0BA/
Uambojy5XGlHg/yXzRIktpdODgbuEm3u+KRN6bCpEDislgL3GlE9mOZTCxbvTGC/aE6nAxfaJDsY
WQojcyoedp4Q8V9kfRALacaNmiQ90CadSt77MXPc1OXLexVSzva8pU2g6kX6yJYJrpgvB/k5sEbE
XL6efwosetuZfyO2VNjKGQnOHUiHOY3tUX8pfZa4eojh9qT1FXxEEUT0ceaBLeH3GyhecR96nGvW
7KtJut47KpEpGWkeCWOMQPhN1Ophwdsxs1T+MsGTbDy3sABSpfZO1/OPluAlfI5paIhDG3KohCYg
BuxzYmprPTNKoYwNkLx7ouu0CM3kc/uvaLAwDbA4wgdndnR3OAqvkj3mtIPgJqSRxfj+wlBEEGEZ
6MGEu02NL2/hrSE9ojj2ah9B8s6nbimYjuycbvxvdlEgbbYEL1vhSEVvY+0uOR7Dsm6tPK3UWuWq
l+3CLji9YixJHeDzLUqH8pzWADtgBeYmmavnw0TcPsERGHm9IgscYwI0PvTlLaYkZ9MNIfGHn2Im
vrBhKTz8hV96emchC8hw9BmZ9QjC69IL6tl1VvF4Sm1c3xDu1NGj0yCv4npboiI/ub8gGnixAc95
uKGmBOUm2e2qAftOIDTn9LFV/bfYpuXqepKOGXjjILKGIKhcrdzILxnoKChlccMGAriK03rGAGSg
VyS40lMeLr52L96TBJIrZwX+0jgfJ/F0ztnEpldKQKa5+ZuLBQoCOOsAOeGE+f2fsvA4wPHHx2ll
WiIp4A8rOQpTk+/g83alixtne4ERmW/vwB8jC3QYWHK6IjnD7aLGKLZpC+zQeE0pxIA5DGoCN0DY
mUiO9sM6lH830qNMAEJRfpimUxiwvorzN7Ne9quI5T+z0LFW0E9SmxJsG2jXXeBB4FSkHc0RhhwS
FRVhCDCrmER8g2+gnDJ2Ma4BBRi0UHFiNahOvHoCDmZl6uOqgSdBC7SQKQxKY0sP3SKSEJfbU4ct
8UDU8PpxxGnxoXktSpX6NJUEwAv0d7nFZhvizxyFXmLmIWC4LmwCNDEypvFfApdEZTTL4aHFa63a
qfLHxJljY4yFPJ3QRE81RewnDJrLoyI4EQyEvxmZWtfaxLRsk7K7ZVWUOG5zfQoSKiuEhXa37qXF
Sa/mWPEgTXeGbSYA/QTFeQXYaDUPwQrax3w9w1+hVV+IoJnmBHJ0r7o9ADBdSTem0SS+aceok52u
4DFnEkkiBO7ZUDunXrsnWXTwq2JB7at6kyI8uZnbTBjwiRR87dhEv0L1Jk1QPV8PvQbjM5Bj341L
/SiAlsUc+mXraWFuvdC6C12eEXdy3t+U3Z6imA/8e6q7WkRieadZ9idjyhycjiFRJiTttem5pjwX
8JuJahzB530eR8HEyZF0xcXtOqpSonWsi0dnMXnG4p9upd3wA5YfMMSMvV540nHvMMTtcx48RNhk
6QfLIwPmGG7B95udqDQjfne4fWo4kkU9zAcZ7z8IFbscmA0q2nUMTjrjd4N6eI1bEn8rjOTQupGw
d2YgjoFE2pdCcQc2tjmPYHKit6adz1hglvE1wm2IeRpS35aTzNR111qSlKO1Zku9galBo5seckaF
EnD+k7bYXtyUrNIqKfBvQ0SPE9xnoUQq1Av8M5aUZh8GRrsDxWuakMfdvC0IgeJc5O+TLF9ed/+M
Cq139GitNnnL7dVj12roD8oHnLMrX8c28va9KYrBxxauc/FZLy+n5xzR5lRA52jpLCEJP2yC418R
TSONAuJwkVeSIPkAzLSSzooujLnLXtTH8lh/ZRUVvt2uG17xNmvGJ9/bztSnwun7SFPPGXHWEypO
azxCXk6pMlnI2WOm7apVTKeVrXphxv6JuAF+ArgeoiUNH35N6mBEOXfocvyv7Aya5+lXZADWVOcg
qWkesAJh9ADwbR/eEQKjAjW1yjEVwsfWP4OgNKiO/d+7qJpI+0YhDdVfkof4mLmiAUtP+8Obfcx1
TbXKpmp1V+ugMq/FHCSbIKCQca6Ozl4kLFWIOqSKHQzKc4CCdv32ZHNmrKtn6iqmEh8VVgOcS1W2
Jfmd+6PWHQF0GVuYX9UN62PfD6nVknoiBV+8BloCed5VdmqXhiCID5ZOHd6gYUqiV/oC7Cz3+M0m
LyfitIeejOrSRIoFiJVOC7Lpc+Iz+UR2gq3m9Av9Zu/HUd+rPrnooouUURpjbT4jYYgYk/7aNIST
iLE1x9qBJlf2/1vjdGa22fk3CK+5VDnO1cZt35i/Zox1V6v8XZdSB+99fRtRE+z0p8d+wOXAEN0G
Oc5T0sqbsAQvmWXWj/dMZqoVcykdoJWWiouRwKvhEi5qgNaR8PdZ+VVCj3IrYua43PYSYsJFq7qc
2eBuLBfHkMp3YsC9gdP42kjoxJ5+E/PAyL9tP0KmBoTuZbdwKHbfxpAzc8b6+nTQsC8ojTTpXnwo
dMO4Hm+tHsImUfqm9ynGsII7lzoLJN5Xu9ssp51ME04kcxdCpdc/M498e+1hKgSpVnQ1Ni9iWYtF
xtV2vb8stAblZ+FQCTBg9UUjZ2KMXMmb0LDP426LFVCZcNh/UbhpnDSxUv/WfaFTf0tooKnHAVAZ
3cvdAhoAMOEEdh9SXdqixFH9OOWe2WHlOJMVavPyFAVhU3JOMvBVT+thff1dvRB97sPbgZmHoh6+
BeSLCGYfSnsqsNR6s2ff1+lDZX99BXp7bAkA6RTXPlooMzsabeKi3nx5g1ifzFI135zuHeg1JjOy
U/1e5fzkUiWylgdd3yUok5B9aRMW+AuV4RttkozYjYxn9YQoYQShgoerwm1p1Xez44xND2eYHeWl
cQPW38HfwX7kzkEjGWSOSveUBWa0ta/7jr2BrUJ8I42J/Dfn6mv2jRmA3pBGqI1IStwuw7CePJt5
sSKANLVCiZcd/IInqZd0wjhKix/6PNhKcBtTHE21WgU2LuXMdwS8tRRFzjaqgbmhk94aAL5B8Zto
3wfZw7ayVPKG/7Dj3Jo0Gba8cin5LA28Fqbiu5TLCdv7ztEwHZ+nIHXN0MS2rRJTTohs54rq5x+f
zXlmfvuxZXW4hfLy5G7wTV1R2EHvKHsrHCszoUpee+HXxNZaxcuj3JCAYvb30/qmc1CDIGo9f/KN
4yJ9RZL78Mb9Y2LicdowzYs+AGI9tXWfVBp4G0CHLA3Zmc4akBdMWLtE/fd+zl+uoD0kR03cOJC3
9u3dhZ994BQ2hU0909+hDcaHfuF4fRF6M/nSjUcZOeHkExPIZc8JpV5/ipoP1uGdPQybvi7964wo
vDcVMkUFWgIT9fnAqPSp/vwMk8WIDQFLjSWU3buBum8rhPbTmkLnQoY2TRun0ChyaK4A5vOCEAEm
pj5Tb6PhjBtv4L9DQXfa/nFzD2pgWOWEdLh8vFoLZSOFLXTVnb02TWSkhp8GbLZTmHVLfX3C3nZ2
NDPqDfsXDPgH68iIhyOVXcJAOVsXrk33IlTQQx4yPQjCHBLEIJQTB/niZOOHaPt5QZ74i42NcBTW
CoPKlOmKZ5uTSxHE9aFzVTnW9dFPq6tuSH45AY7/68LbTLOfzXOV0jj9ZTS9XSv9MiZgH9k1mqIu
926pu3wVsmfu+wT2eaW3YlZBlR9928UHXuXGaZ8X3cDfUBR/LIezXFOyCJ8BjA5GB9P5yDVn8Hsd
NoQCnoUB91E45lsJJ2fDK1QZOh0sCz+54bMwwPw4g+Q/1YUrZzt/Iw5MpCfjzIq6jbZMtofSNAg4
8zekvNxsx213YJsyH2o0zoJWp7WN3yjWwWradwfpt5arAAkB9Zjp3kIYAQ8t7nh/OhJt4rQ9I7VL
OXibER433d26WvnZLv6ANGMeysMbAUujOFsGtTf9hIVzpdenpYZCUmnFCdABAFGfOEgGrhbj6tkg
N1LU9NVa1JJSdhQFKETKNQW/kkHUjISE2mhWia0WxwwZ400bO1l8YyvKzhDH2Npn0XEOogGOyEkZ
utztqGQSNsvErTIH8EVrJpAqppkdFidmekacsp2EQsJATydnwCMxgp9Z2sbfVZxg30FFyPqFpJBf
MjGxJR7bmn76lB1uWRTc+gn3khnWyERQG7f+D9keR+6t3yjfpn0lsHnqvqSyZHogo0ZUtCJ6AQk3
S9Bs0lGxKa4niYuHq6j5tkdDOmN/RZev+cEaaO2u4At/tPNeBm7VM0b4WXR3d3wKdJY1GGghecfI
bHl+HZAX6+eU8Jjx0+0cgi06lQOsl8hL8zQc1JFqG66S4WCZO5d8JtaxEt1G5XO68exhfIOOcJIi
8viVFM+H4xvOKTGJM/xZbCnFckt/fqMa/8CfFlb7Og72nfA6KxyJmtFH2B1FK0PGFEN6007la1eI
QVquujagPfCSvOalfo/gFsQ+QTHOvUMHPrq1rGevwaTSNW6963MjbL1lEAkJfS3cksc1OKuS1lfN
Our24BD07NSxo7FS4o2LV8ULr2rPTFQfG9LlHahRISN0LYA45t2CLwVaiOdmk86HpXrZeaUtIqYO
Av/ZJ5Nf/odGiReWt20DjSBt4AjHi3IpzdqROPwFnt4fRQz4B5yEbWIssUoyZsu6/gKmMgRHEl8h
j1OumpAK16+kJNiOBW+xokLoE+OA4T8eGOeGAsFD1n5xlKjoNXqezu7SjP6L5+403Ukc4IMnLpy2
FRoKDxNC5oJPSGxOX080xE5//SANRFOZdDPm9yDFrQ4A70pNwO77H5uhyYFa1wf1PhkALDHcJqMN
sIhLtajUr0tpH7dSiT8RmZ/mf0BXIEiitkSyQf792JtRtoSno/ex++D+KGLdMipYAWRRlFDWsnJA
za25FbHzd/gDXzL4poW1T6t2SAvD4zeaFBExxbKvCQSrna9QCS2b9wSPRXCKuH7R1JYqgQiyENIB
/N0Jxu+xJueWxAggibH482E6nIStd2jjExrnKdITdzbYFyDdSMcTXobU3eqdtTW8w2JMQ/ihNWtM
AaV82VnG0Z4kRrD8FyUYBNEj0O4bkQ2EVQH9uh8Nx4Vz4uEKPZonR9vjOVzEAFb7J1CMMJl1buC4
xUWN9HQHZtR+c9sPWe7JzMhOF30uv250J72L5t6BhHkfpJ709FxwQVzRYiVGLX7zko0MjtBQzWKh
tD1v0SH2VhXPywnUlDqwAj5WVjTRo5+dcCTe8TFZSdEONyz59q6+pG4R+LIqJAF5TUN2DpezhBck
c/QejLM/avQjrbZNVLSxRrfrHAAmHURSq83ALXlZ/Wa7JMlauKfTBLjcU35gP+VWGhMsrXlxfC9r
byUlZ+x7mKPsP9njMfpt/LPHoDpI4COBcDFS1LAnykEh1GfugTaIyIYGs4Tf1F0s5tK5U/L1nlv8
hq4cHF1t/CLjCx8w16o8XXIouWy/U65iaJoXx925C8kKwQ468lYi7p+3mgevrl2g1PCPETR99yDL
tVAPUuHE6D1/7hoJz6wByhUx+WYCRhMuB7enRFuoHos1wBQfpOjse9ypW1i/WpATvG49lFK+E9ey
BoTyMrSOPj/6Cat/sf+3CxYbb+uuyV2VxCceCsnNFa8NO8Ek4Jdn0YmvAlz7mIfnz/Pe7WCHZKDb
YpuM/U9fI6RZi9CfXm3DufwDGQKNnCSlH+sZjAmyvpuTq0xG384dTrYh3LzQWys67NbYGNYO5qTN
R8TlHFYstb7au+sspvMOad/TMNZqs3hjWyfbhL9b8/DL715//69MIHwd4V6JdDHJzwEQRMSS0Au0
abCD4Wy9mMt8oDeKRt886seM8LAg4mA8FwTYFe87Gdv4YZITXTk7M9Omfas41Fyw2lj1W3n/yAqa
hI7iEetNvbbdJaawuvTHe9SYnj8R/5K8wyYa4APLLOda1McJ9MK5xN+zQlKHgJhP1XcZG+k5b6HF
huCx9l7VLIXjPYMbBMyQGI1Z1MB0cg/nV2wcYrM/olMWS7Zj0yq+n6SqQNvItKQ42b32KD+i39C2
ryRiwR1VXjUg2DOZp8vsZuOX68XXPJ0aOJTpqTNHQBI6qdpNCtmOlnhfuO02HdAMlsPqs9ifMynG
B/XAFwG367hWy8GMQ1vytEif9nazHrF/szL+aMz+K7RMNbfSc9T4ceXCEtD16qcE48SlVAKngRyc
JKDBSVtyFZ966hQzO7msJau46Wu+yIxP8BNiQQI2ho8D293Zv1cGYCnXSY7Shyyeu/VLfAIPGiea
ZWtcVrsVb3nZgXV1iSThfbaFkJjnF+WUjos3yUtCShgMN5CXhF95T6AtTbp8Tva2EKfbIMZzyuu0
EF04Y6VRacBmnqQpwoSaIfHd7UJIazR4IK4FdVkuxqOcUXu2RldrIGfZ9ISTExPzJYI/ylCCBong
F5a531tN3xR+aMacvTX5SA+OJgF67BgjAAursYzPRMcXw/54BVrQMfAJ/1z33S0aHebqsBaDyfCc
VNmsDFYvZPclGkCujUEu1Iz6d89kHWhwnNppWL0Y2C0vaL+xn2k1GrDnlw853Mt71L7seEnhyo0N
fkw/OfgVU8pa5cB0LcT2TtxE04yIVffoPiuqHFo+O6sOnjjoRta1GNkmXpSe8dmbh1y4+zNboOhb
w+HXN8u/qNOnzV9oHkY/EcUeYtArjWqytaZFthMaUdSZYXuAPwnEwOg/TLou5ZZCn4UkIp7XfoGm
UhWQXvU/acwdST+AXIhK2OWu55DPiDXPGhFyAh7AY0CwB3DLHfT0Q2a8pd+BcrTkLxM4SCIyCfcu
6A8+bX65U5eS4U1mVgXAKVcdRDRRljo1Nwrfys2T8LO8Xj2E5/DW/M2GZGUh3xNLNN06fkW9ewVu
CJ3kkWGiLKzB3JUGN+KLEHm5/lV309EvKWtJDrF0V7H7kAY3q9YbvIzUksiCguVMjI6kt706qxMs
QqPpxSN48cEw99WDIKRGwA7uyuACFIMC6JZLl/nTi3czEelkEoJdIpSkOnbUDWhB3JPb4IRlbOhQ
w3IzN1Mb8M+l9CaDQfrpIoysV2ld09Shmd834nNZtHUpl0WACxkla55052X68rswcvaTVGp8rke5
Q1rTtvkoPu2MPCCQJm1SHaK8HsAuU8Fkz4jHBLCq2IEbQgh/TywIp9a0HcwYZAgxVZSBptIlinve
UQA2PRHmGH/UIcOCEXYtEl6Av7+Q0/6ahIGBBAF8fAzS4W7tGR0pvEi7gVuQrovWT0SuBtZ7OHDl
VCOGqDGtJdrzXiZeNTkytK/do9elHxE2Rle71SArNavnkodzov21eUK4HY4NfbHOsXFgBlwlLlOo
/HrT+v1BBW22Dl+9oM5V0XHAcmszMNPw0NuKLECSlBNns7vXk84azDYb9AzCQdI82BAR9/BS33hj
lClY4XxobZlE+ds9AlilLBDCu/6dRvqtB4KXSKHu3QlNJnUjty7rWXDTO23U52PYN/zRyHCsS74K
Vc/0LzaepEs2SmTGTbRyRJ5yl9bhh9MjYDPhaH2H251AK4bqGyH1Jn1MFaxjrGF1eTuVUw1eKgyg
Rdi1+Nm1GKgNU2Z0DK60bb1j84YFhwOyPxE4p8tXZi16XgWuA5IfuT7Ojv/vAoaMYWLovmnOmkBE
axBQKQpuSFAsXPF+YH1OD/dZgKTDZR7dFSsdtRj6wkUu8ed7b/atSnpnrdCaH3ocNXFzU6CVy4jR
FfT4QnNZXZ53lWNotqP7YXG92ZsvOKJ0QZMzCfKmRqSJMkv+t7fnZurOxhWMZqYd1rrkNCsyzJx8
pvjFftCFzB25+LWZ+5zJ/XsdB3N8R39MTFdS1/4TJnEk+cf/DgfI0tqpiN2BSM0PVfAFsedOyFvB
WEj4T3T93GR8ghd1HajAKwoADLbhr1mDZOcfGJ6JtguTzW6kZzNe7mBWc4xv0AvU2vJZgYRviMla
uUnXk0Vff0z5SxFmMejPwlW966JvsmWnUQrMoKi6DOUJfqxT8w72I7qmbu1q6xs08IcKSWEki6o+
7sZ+owl4G9zxSqDSMqDV3W5sVK8C/MD1m8M+EnQTP6bOurdJfOu+zmn981meM+k8hZ8bvsWx45rd
V8dWv6MPCYP9EP3DzU/GFAmoEGD3XbDuSKwkyarapGj67+5Z+zxYzE6HbGUbn11FCTdePKTSZud3
gsZiR7hrU66sMSCNfOAVsy5ICgOMskhOcPI1fTBeDFSUjJWAZiTrz0/vzwQxo8FaMSaayOtd7DfQ
AVKWkouO2sNlatLeq6d0fhWjPKToqTQ1bDNfiaSe3aU/O9wRFp1X0qget/S/RjrN1Sa+9rM/Eg6j
STJdbCeJw9VxGLDVD4Jmc+tVs0KdGoppYtu8/2KCLa59dj6raZx/8aOaL4kBeApssXr36SG2Wuy4
66T9TYEZTo+OGNZJWAhbxvitVEKNyxh87FJAPUzoinO3Xoe3zMYiWEu846GD01dwCqxXrOF8fKec
rhQ7rRG2QEHEV2Et3n1my2elOXBppyfuxGK+iccuSXG53YxADT/0VILLW96RORLX/YvfURiDVr+6
1MN++pMjH4IR7bZW2BxlUW23QrWBA/CFPxVqV5vEpR1/y3sqSYkCXbr7tMhWdirpGwUCNPrXRh+c
ZhscFeqaL0Gy/ydgkP/RkzTbkFXnn/ou84kpBq171DpH4pSkUHYWmSSDCZAXLwmNyYvvqU/vQbdU
gWhjkHylfWEmgNPZJU8nLh/uY9UFBoV26fkTjJjEddteEshH/3Q2lIZIaGHgXic/SetarSDxuXAb
Hc7ekDWd/L77TlBBet1vRpjeO2xDa0PKtK2/v/6K4vewBeyV2cy3umn0ELxMlch2/B9OMe1DGq8w
25+22hWjmzjBJO9I3DVaxAytYk3owpEA+CDMHSFd9juUVhmbJYXScyrGjL40g9BuAgQuTOFKlsjU
v26vG0tzxtZeJMv166O69ztvFAOldM/2bCbMV7RGOCuy3L939AeEE2kZ8wvbUqe6CF3GbgbjbtIQ
KzdPrlVmFOd+xDeqW0wNC+ag9FWQnWTl3zEgddlPSf7qxVaspA9U8X2+R0IeZjAQ9k0nXIJqzLXg
AuhRM6sa/ugq2r6EIGOl+dFWY+djk41m1rsYyLjpELyls0tDXojFvGi+Zg6EhFjHJ1eJXEu7gmpM
ZjqyTXWhumKQkBCr4k0HqY1PU4EzcSYnP2ehTZ/fe71x/qbxps9otks92LVWcaJBaHzXsbgnnMZI
hVSkaeov6qRZszr2uhjvJp+P41HFUUDybXWCmhknGFNnIn5YbJum3GdUqHV8glxD8p0pVq7FtV07
83bbHwAmcxdYuMyhi40iCs/8fVoX8hhRkrtQD117mpaMSnsGqPzYz1heAaYlCyrzzupL9AHyicwQ
uCCtV1O2FNftFCHIGEXWa+ojeaHDiyx7IFqdjB7TZkxooZ5jZV6YhgNpDnLSBptK/ZWd2bDZlqGx
m7Qna1ndBY537+IpEyZXznTrIfABZ8R7RIEGUVIemCLbRuwHWdo2cvb+nBlUhipu57B5/iTgnTUZ
pGAFJT8h8jM0pwAvebvzuRxsHaHShJVLQ7th4JoKV4qzMWndusM1KjXxhuR1+ovaeY9r0gJ5wY75
gRH7lD4jzR5jfXQU6ENjADnWOuSIIrO/kWbR/KmkIAaASq85SXpHuOUesqN3DSR/FFrkIDFbecAZ
4N/F7PRIk9aCNJzZ+nxd5X1d9O0xS5wJYJfxnRrfY7SuSreiSdUFecrhHhe5xBdAivNDSWL704jc
U/uMrxMrdLltxjuJOMezH9VY2zHG3eFPyKcVjBY2bu9zVXinbrJYVdwLYiPBYTZpp/OiH4l8ew+L
gA/WZewjlrYu6FT/994l0G/JqTV+RA/bdHl5Q0mMCdUKdx5+cDniA2bME4jl8g9s4/BrwzVmGO1Z
cmnLPYZ0/0LgQxw5/rmI2I7UttaL+4F9mhanffzt4e5FkMSEsytNjf4A7Dq4OZdD+a4aOUtY2be7
563rENW2X2ASq4IMmkpHvErOURtu3vgQaHTzrIuJSRWjJZK6ld3cJi4RY4uVrHjJq6d9X6aVDqXc
aFy1x4dHokygv2u1aPWRtqO+lECXGT/nPT+DclXIg1VQpnLjd6xPn1YJsk6EmZLzLHwU6VB+B0B6
aHl05KqwxNKm4d7OHmd4a4qtBTF8kSH29y+I7JJaDfaVH9fKFVrRJ1ypSrwKNdtq13FZTZDee3+X
V0dgOSY4ZchrkXC5QEYv/OTGniCFSToX2rNbpgH77plxmQENI5X/zzfvXY3Aj4ts9Ij/hz6RKgnj
Y+WP3XlDc55FXakQlYov4b0FtFngY9FvXYEuFSyl4lzVo4CcR13LvIwBAAC7pWUuOG+Vy2kfFc1d
6nd0tXyA6sQFMAX0JKMvazuo4+QQvMTMUECsZ7EoNjkD7v4E7Xc56CugWF93Vk6OESCi/YMINI5q
B00FetN+zoIUvzRZW+f8zSZ6XZQQ2pwMULRuLHAH6Hf9GxhmOenmuLwGnWLu0kVXn7PmnzWLmmAi
DgKvShXg0MFlYfJXOj5kzc62UeLwgNiHrEXnYkcDDjJEFUVOr2peyWG0uxE5TBuiZ5hHGucSM6+I
fsewYmtAmJcxxLeQJzG0FyPq9zSaWwC7CGdL/CGmeLLB5qEPU4lGDTLdbB1ATiYc6Hj7lnc6/XhJ
sI0Ir1OA6rnQf7mO9H7HyhzpX1swx0US7UESx0lT4zSEWQDUUpYwtMjxQJ9mHgaQmeHvaN11Oicm
rzfA4+a2FuL5qv2UR7RaStO9iX+Cgovp+TT26ScGyn0iFO5ij964xeMQrSM1qVzsIBTHzabxnxwe
V3czn9expKJhpRdnf6/gJq61UN7iYu6NHjuQuJTwtBK/KbgnNCZl6SWZ5tEAE8Ag4uyGD9MbSJMG
jbaL0a3ErDF7nKvMgK7jQ3rioMYfL/Pt4dCwtNmB/5ZRRRNsNHY6c5Dmf7mqt2cymtSm+KR5AlsI
umQhbAyaN2fldnkCzkADQGmk2WCRgZbv6Z+EN2+rkdMTIrT77qwardD4WHAEAs42lsZOLfE6HLAw
eT6pct1aw8rZ9RsLpr8O9AgSFT24ZDDDpgBEvfeymHGu3uEIG5LdCgeWoJU4QBEnbBfR7bPLJca/
1nbV7/FIFAWhUN9zREOxGd8JKd8Y7ZbanwYaxksHf4OWi4GhnesVdgs95hgX/YJAVRBKp674Adev
cwIHDxYv0w7swcVdBDeLVWO+wGYh+yp4loTHTtToGlYu8U58SSSnKSe/XVrSoS9qABqH3NHfRu/g
OcfTpspW2l50h8RRjBPeb4tphogpdCdVq4rPCqSfKorUySMKrsywepCtZW8+hRPXG2hcnKkd89XB
TJEDDMSXNhGkjAEFopMqVGFLh8y7q8yuPkyRWzl1VLzEZETZenFlIzxG9zTPQrxXqkfKqFmc0B/e
rFQ6dQ02YeI0MHcBfg/qh7vXx4OT/Xr465pRu+LhL2V40gpgnnQKMHGT5Q3C+Er6J8/Evr+u5iry
NknS26fejFUaTuHNOguiNyaRF3ZVhCejeOJwfdYV3w6wQn+oQwa+n8qdiHRGhhLdOYvStdc2FbjL
98OhO8tbwJ57dxsWZc+syWgKFYm0Z+r751c+Rl2hE9RDVm6q8d4vt7fHIhpZk3fwotNkX79EOhl4
MixZo0xYc2XOGHBIU1+jpT9eng/IHQnzjGCnLbPZKjULTEmfYeXEKOPfamkGxpospyCMiiev/njI
zvrb8Rm75AyRcYU7Ua7Xxt6TXkAbamq9UPtIOwj3MmFmjh1NUaZ1gkXEdH1xTZtXtDtR14DYHY1J
yH/IdHx8YbkA4L2VTfdG+Q+xaJfHg1Mmk6ZZ+klmX3EkBXtX2XIgNaghky+mWebYnnmkf3AZKysC
JwJYM9HCRTgxSfbDPxTI+ZcRcF54HMZdE0vd6bXvQitGMDXx1vkT2wXLvxRqhFpAeQt6AmqPJe08
3VDyRJyjYdXEu24+wEMqGOOpKHHc2/bIg3rD/LJbkZOQImzwbxGz96rkhtxe10k7ht1AWMoVJpOX
ub++bMhjClWOkjzKzGDAntOqBQAjHDRI0N+E8DjvxgcDa68iWMDcTn53Yr2YSFV0st0CUFgeV3K5
coi+Ut01EdLjQW5DIYxUiYdBhYNd9ifPqdqRnw1mE7lpC8+koCwKzncM88P8gfRaL6pkHopQHhsT
k/cgLLJYhPxt9WlbmIUF332AnPW/PD4nw8xXt3QkRgMf4yp3RXzpfIBq2W47F9EerBY4FlPY7OQA
QehlzG8Pq3NujXwhf2soKsnS1xtO8ThCKEdid+pntcoS92eVwYIYW0sRrwICwh82UnW4VwwTvFB/
DF6znC2GTIYUaNxExLDInCCwbCWM+QHBDILZa6SLZfrYxYYUAwfPhCVuXRL82nFo5youl0cODS/3
A9YPf9L82/M1hSDr4F//H0h3z48B/3Gb8zxwcUJUGQczUaF1Yb/BW83z3liCbHUHDrTuj0eISDyV
mk/olF5sr1gYSvKD0wKk2DGLprPeaWdDO/OuGs8wgKvB5iiwh6awtxP1vlnjjhi4YQ15Hqohg6aF
TAqHCNjVlfN+seR16Iv2aib9LdtuC5tJix1i9hdZPPoKVWgKdaUgku9Aqoh6bzbIAKgCIdlTijAO
IQn/2lAjgi3Uus4QJe8R8C2rr2i4P4bA87Yg6pSOlDGmf9CW72rylW522kvbDih7I0E0/ZsgqSyD
aruIU1XkIelYYzPeQPCfYaPSvaz0mT7WBLNWt39n7o1E3iTmPb35odbmLT93buGPpakFm9o/wOTs
EQ5vdRDBnv5OsW6Og9N/wpSFUHgn6oBspPDAhzFWpEVigciXoikWUrInXjsrSNmiNrW5OiQ2O0Lo
6NQCHYEipCkmRacUXogGWdGunLmxzW++xnf5TKf9WMBvkOr9cOp6aoJW7GuPbshQX0nBPDxOA2nz
h6DiKNxBMqtPq4wF0J0wiwWicAD5/hqgx4pTjNIIytqfTJBGC42AE3NW62sP9Tu1U13mXAYvP5kx
ohNgkxmfbJKwbqip9Egp8NOhJXq1Z6cnYp1tY0/6gVtUEpI6RfYD7L+U2YDslm6j+s/RJbldpbTS
r+mj4QpDvj/Z+dFYFBtUuhn1cU7dMZkql5SN/5rAXlx95nYKSnX590cl6FHsG9xZ524Tn/5flQDl
dL2sBfUhoeqUL4LHgnq3RwuguWlAidTT0QYDZ/wOxWtZhNnU/ecGR8p+675ZY1BZaEFrKZ6RbCZr
E6gZ17T44T1Pp4m0DVf3481ZKXqYV117UDa+enldf1B2NMDHIBULfeqKVf57eirf7wl+8xV9Etci
DOUeSZP/h2RezsP6kuNSPm87RpY9go68pVeCvQ9KbPVrpqfUxbICYCm0krvY96TRAa/vFs2thrYz
S7tFQpuOgZ4qV9zu+B4qS+MBo9WuNYlL038kXdFvKdWJAv3aUZdrmTLJb2vOzZq3zZeEozDObzd+
pW+QtVo54r31NsMSo/dZ4YCSZChstKQ7Pfzc3+gN9gyrXV32OmHJxEIOCZvNBL0MCHum/xB8YJid
7IdV5hSXtn6096KLDjQP9URhSpzot881fwrFXoi3yabWr/m/EMbLfntj2veRenxY2uTxoHhi8a1G
70QrWxxJjbODrXnQMX4RfmUx4WUDGWPpbhE20qaGFe1MZakTTSoXIYp6OgxmL/Jf0Qk9tfGpFzro
TcYjImvoK7FJBV8lniJ//sMSLTejBWp0x3bhnJbG0s0t2AD1vMePp3js9n5hCGXQol4RrwvzwBNJ
fkCG2I7emllNr1jMrVFiJzg8cU/BI1XCPyvPp4G48DdeMTEnMQOJJbIiEAWhUbZxvwnPq7JvZtAU
igjNBSpTVHAYWbEbiMhjVHUbGv4L7bw4uC5DHQWiyTZ50l8m9Y0i8feCLZWabCQq/mNPExtlDy97
fM0IhP5KHGMTuedExouTew23hkQTxiwiA3aSoK1WQZF5BEdd2jiDNp4EiBgJzTcQAimgng1CW6f6
6wMZY3H2kyBmEtFSC7SZvu7BjFmtUgJivAN4L0cdx2ncqspyRFwYuK2u9+kkmCJuX2N1LazGEYj1
CUvTSPKiwhZQ2TTQJ6F+h1orm2YIcbbtUZEmh12Q+1rxsXemcrF3EhJoGZ0hEgEk+PPRjAbsE9Rh
Uc0jjFNsxeapGku8EtiNzVIhDRhu0+xQrf5dbGePES+dX9qPntRvDWL/OlHpHbT4XpsQpA6Y2YUP
37x9ao8lr08EHWeYSu8PtH4Vjgw+kZD2xmstgX4a3ou0RpWDKEidVIyHJsgNMTbdPtreGfcx51Bg
dmgPWKpBjlRTXyAVPgXA35ao6mbnyz9k3vnPSMJrGTivsM92yXX4fG4N8H19BXxwzXIU3BfrTH5E
35v5dQxYXWng6FkvjY4iKLm3E3b8MS1HLDz6HtD5RGXxeCLmIRqdj5Jex6p8cSfVe6ejD6igl/sa
hzjW/QCVFdrciV5KVRxaRtq4OuNIzZe42wwOcQPWGbpZsrE/YD8MdMN4w8msjYqdyfMgMYM3xbf5
8dr9vAQZpAOUNDs2dZAKH81/xnltIewDPDLgjrjD/vNNrfdCRy3sfuMwkzamkGOM5WulQus4zcH1
emfQ4NzlY3GplSTgQdfsFRSmHemOUe3MRcCgMyhwmlUnwJxbflrxP33hxxE0ickkQbi7HJUzT4wU
QqqWGGGLgO6Sss2WS8Rq1S3oNKi/zQqTPZMbsSAB0GBXAN92lM72s3/wVWTRKiScvi2Lmb0U1zoi
W9sIw1zU93HmLC5KBF7k8XD3gcrUv37g8xSlAIReZt9wZtP/Ut65jpv1YZVKETRDIMD5Agk1LnkV
mtml8JzoH6AMHqSQg6N8rBiGDMNjbHBLAwEHxar5B12l+BkolGwFB8ALgadyPwwqhVneazug7lz+
HbfESvJ9dnM3a51kP7LtJpNcBqnSf8Fs6hTB/MxW3O7lEer0e/1QuSLicy2dTBiZwB15fEepQXRY
YHHAKGXpT1KvCWO9ZqgrFqIuCadYj+YnjhKSqnrk814yB0SaR53UlFFdMmuzvpBtYPU+QFpmXu8C
DpNhWgFpwafUD0xvnEz6geLOuDRr8bB3ucD3GWEi34HwDmw0i8FCMsmLbKPbpiX392ffg3IkMgyM
qL3Ahuv9249Hpgu1OO8yPU3E6CeJXc3+ZQ4p5kSgGlv1Q91LT5Yo1NGnB6p/StAtvJoUYLCerKZP
udoDSbSK8MgMV8VuzAinaxIY2v2jmGbx+rh4Ec1DmEirAJgDaVqWKJNQxdL1nDZ4hB9GRBUCHsXl
6+PSSe+CkRA+AnnPOAzwCuoiF+CWMjqeSnA++FaB73L9QQvVLDvOfpvuCqquo+7bmB2xeZneUJ3z
RmD4jbpJ545T1xKn7sfq3WOCkWHU+wrD20g3pLRiBQlQnMiLRPqCU8cXtWsV5J/r54rptWnoVMkR
SDlSCTJJZZUYlWXw0XsmKphQ2oGqaYVb5lz/S1lAiUirTWG+9mqT8dTeyKA9snSoq9gpZOh5JXxZ
iVYjAQA/4Xe1NN1jJR9W/Jq/Ld0WMI5iqi8j3mixNJ9SttwXrockNQl3RlA0GUDdeAm+bnqOMfyb
yF88gWyq8sdZgKHXRnJbGqEo+7Vjq1+EuoJAIXRZHi1O1KtJyze2J0AdsOURixy/KZrjYJp1EOIo
aQjVCurn/bPgqZjbT+lL4KoUEjBr4w99LztCL+04gF2Gbp/uf1Ny6ccSNw/iGnl0PKKNyDf/jJAE
S3855cIx3kPRDJW+i4d7T+yeycW3VWhH6iD60tE2dMeenKPu8bVIVhgxX2r0MvWvLSZBo5HASuU9
SR/EK/DKTvsHs9gEcJ7VGeKoWx5lDCNAiOjAXya6JKxcg4ma+FEqhl3PLgsELJ5zrT578hVYJS7r
0OLFAh42wqNnSWacT7YVM1AU2C9geGPFUTfEIEiRLQL64RBBauAkqXJ1UucJ6R6NzGXzmd/OcL5x
xkThvhDWpTFgsfNxiLaaj4F3dLUktRJ07w46FDWRxcZK9bpwBKUuNmNF+AAozp+X2z8nEyxZwsZk
B24tvdayZDx4Np168skFnwNGGqweBHtbPYjOSOL91+QuD1DTbrPd3XKcofvCDhQy49huy45JSy5f
OGVuNpzsVVPR+kVATtjTc/GqBu8MpT6onoXfRTpYQyv1R+b2ng9FoSzl51hDcXMao+Bf4gtBwOS2
PkJSUXTjqESU7LzfQI2V6YAEnSoqpSi19z9Svlher9hE05xpV7GIdfQEKEmE7eIyISkOSIKF8Qna
c7QJDnyzlpjR+h421GtxF4Z7Rtv9G/eHy6HVE8fnHH2uzvyugC2GzBN2S4YcZ9IqMDH4NE07YHbt
rJSDQORSzj1vgaIFlhkYxYL9MZq34UYC1CO+suYe6E5QRqGmj6OCb7cjch5az4V5aGrZtCwA+xMn
Id/OhFitPmqE0pAXDp6/wdAO4S2oYfQiQ8cM5Cos6JVXn9C81Xxbk/bqu9TgjW2YYwXjSKjBmrBS
3BTXs0ICrwCSxhszcCKuz/y/NcuD4dp4h1e52/QuMc0ad2LmeRwF8PLQ3gc8jrqTE4fLrD66+oPV
M9wS8BEPk/NMhLePoGzZPDvQZFNsAPVg4OrUMC4rLmXo813e1/uLS/u9q2QGUMM/pwaykmD6INLn
M6YAtlWL+aKkPsaYzT3x+sU5ZTifZyMj2MG1bMP3ueNpWG2NhsNArPm385Br2ofZjMrBzXRapeff
6xLJd7eOCuhwoj86ZFz69fBhO3cdAsNe+8jirZq4/zkCkZBIbMNR/p+cqYzn9CTnDtKN30iQ+rXY
JDVU6jq1NWvrVNpxh1IeuIzSs/qaSgwtEFG/NcZ4esi9O2/KTuYtYWBEWcM7n/ygHvUm56fat1/d
MV9PSWHmA4NNZGGIMspCZPucoRiaQtTZD1jpso4Ord7SPQedGMrgBbrR9+h6bgkg+g/VXRo8lqfj
HZy27gv1X9H3bAcssmB6EQNSyl6nySnvLf2fE5sx9nEZEpWRurDRPp1uDwiu8B5/VEGBhUCWAYHc
xPh/3GGZSAqwZjjPhfoLdOGZc+o4Y1AbNWKK7f1OKmHPUJ06uoqDg4lv+fa5SKK0UY30tT/aIG8J
gk28cklLSUQv6CVbCbdkQCGCSGblHvjP0KSDOeSoLw0qoh4AWzSLwA2njnIQpzpEeG66KajO8oxB
TW8AwBirAnUlbm+KRgPBN/0Wgygm0mSzqy7A+uzCJwIS7FkPP1iPNE1CmE5I0lXPwXcliA4X+2C6
FekrKeIYCQk6bFwFPQgirXL0HkCK5s6Ga/LzhA2fP/HniFeMLE/NqyNlrTkqNhk6SbaGZdcDzfeU
XGgz9wZmQhJ9mQq3rl571qmB3p8DbxMg86tG94UmqWCMY0l5liWdMm3Wruio7yejBliKOtsCogOs
eTLzRuz53l/tK7GhoPYM9k1/MvmjR41YrFf1pjDuaqQdojZyJMDZVUS3Z167G4jmGXkpEGf6RkvQ
mXt4FBILQEoZQhco2RPHggZaTYNmloCKK2XeQlEwUQOlwEJ1hWmAkdrHao7z+gRHzTZmRLDfi1BI
MB6+Bl6rrjLus6KMFSIMLo390j/ihZw82lRrHDF7rJwkeB6PTA3R1elBvxhPD0R36pKF+UkuoYIV
AtEDcPsvx96Y8+GcZwR8Lcg7Vfu0m9TKq14d8okaT4A154pnx0/GnhbGP5WbP5yM0UOPhMuPx9ml
gnVzMcQLA7JuFzwnm7vVCteRLdKwPiqZr81DTLmjA1RqTfb/Dvhz/Lq6P9CPM/VXl3mP+nFWSwXc
fXtBXJQiRsVclWmEakNExQVuzn0ppNWBKsm+QST/EUUzV33HywKtX1rIG7VcGmG3eAgR5d/v8A9t
HGQjtqEFfShOodgtCerL//uymxCMT0v3559qqIzGbJ8uZqcmJZ6WtNbH4j0Eqa3d58AfJplcDFQ3
643Unm8L3WqWFC9gJU7Lh3vOKyKPBIpOjLAZ76qRa4L/dhFgMG+NagHfUGXdSIjk+h2fIqJUce8b
BAtO29zWx14dH2UtF65PccWlqxzpc4It4FALBCVh6ubr023sguNdZGSWXfOHBnOO/gydki6LdP6u
N9mhfMKTRQtJEUUxb2kcq7FCwsg3LmLYYTsXyAWA3pxYr2iOxA4sbM7FmEGGhfV1eEDupe1sBVyg
o9npSrv5LubttkE1bDfdfXGCPbGa4v9B483C5YY1okhDf36XOuS0ubW1CU5lY4Ydkc3XK+5Puhgb
hH+oI00c905kOWi4FWhh5yc2liRV26Mc8dsdaw1OIMdJFqkNMFKLS9PsKC7qRXBQsypG2vsrAFPH
4AwawLdFY2i+YLqfURXd/UcLJmOGmqTK/1jaUTYWNu0zVawNed9AhJJMwMp4Itjlg04mfkSj9KF5
xnIye0EruLCE+oH2hNqyhTIeGZMtE3a2hBpoW3fFmvVDuErCakxxESH/imfpYp7QH2oIki6jrj/Y
icga+ryXIYmGSWeR5lG8ppKqorGHF4WealJuWkitM1HkVTiXL1PadIAegOodyvo6DFoBkXV8ClO9
X7nyN0n51Nd+91QlrN2mUHTmmgGjQ0gSidOdZY4GBMq/ww1hXcg/CCUZlP7lk4EVNq3mxmv2h7tk
vXNIwmbs4ZI3ezpXlty3UdECYfU6dtrKY57wCLbLfunCrQvNJnWe6rfuCnpLVEga352Phq7cgyEw
IfYaJAXxgyDFgQxOWUJG/MjC7KvFSRN5Djtcah2nhQZTWM6qApevxhTk80x40eg1TKfQRqN99FYy
ZCvL1PgqD/op5LLktGRmEyS+7ZzqnmMHPBYiq+LXOdMuDfoiwc3mWVyfH2Q3PSk+M0JeA2bgLHy+
2ULX0jNMTkgVC9lf6xIkZa5be9qtBxvOAeW27RvuVmzTjbj0k3USWZ0FQqOfvw1G2KSFMpGWtfpx
jy3XgMsarNv1KAkhIv4jKJVFVuLI90LZxMtFBnT5+kNbXklBnbMgArfYqMQ7wXPk28OGtXKJHPZ6
k9huqJZDKtYtHhdcyYaLBrWKGErp1n5NYQCB9i2NZgyipI8jf3zYjHgfEuxhzFxhm+IsEmek1Qy8
3roly17qQR2fpThBhOTkmAqY3lJMn1m59NOT+eLjhmAFHyx3wBW8jScCZyXViW79/G1oX9GHvHN4
/Seii7Kmx1pzuPvU0uIQ+w8oB5DGG7Qt2zyAMhNRk6IWk6nBZPZiRqZlYs/PheinVmUqQuj/xxMW
2NZOkBhJpmi8yFTdKVmuYOtDLV7M78YFWVLXng0YthBrgaQO34kcwF39Csp+lyid5Yh7TfrMnY7L
ti2dzv1KgP/VeKk9QrU0JeF2+C3pIN/fGanhNaUVia78kV6J30yR/fnXzJ6ba+jZiwQQoIWfd1rS
Ma5zEF3XOmoXxCgjnriJPAAf/K0BdjZhL75wGCgHU5Z0hRDHrqaK0nHQZMu77eNpuI6E0YBw/wsy
Yrfe1LueO/g4N8pC6tQRT50oT8fGc0hLYFZRX3IEoQzmoDmZi/64BjdJRlLMKcIoTgmJcbDTjzI6
81Xg5h547cs5Se5f9B1rKqwr+2z/S/rT5W6No9epib8tvyZeCUfzXu85H2sZ3hhBddh4fHSxohRB
uhzS0NQ63w2TJyVqp5pcK7F+wxox2D3xSbUzC13971MS7qyKkOB6L30QRwVDpMVQFYlIvq1NipWm
HyylVU64gvdthtEiKTTuSaUfck++p5BjhTrXVOCvyeSBTxoztWahrItwqE5U7LGaWv6xb2cEHfi6
iKDq3hIE4yIfS/VxqTfNqjIkT5VyB5wGsFoQqM4VZFtr9dN7C1SEcfTEBoc0yJIfM1erZDtfP7AG
cAdummBitt8Psab7TBOXGFoXWywgSz538wB2nlc84Hcdyf3lwIIHQRqIq9Oe2NJAzMkIV2fUOPLM
/N8FRSFeBEHGaxdFrFvEr2w3v/D5mvHmM8Y1ECb5gbYn9NZ+mIneUubv+lygcRbzWPYu81D5gRxU
XByX5JFcPUTLmDC2rA7siPw/xBO0FlCv1m/WEJsjPpThcuuSzOPKEJbG/3+uITnAGD3JpaZB57t8
/s9ca+PXyqk+qg69PbTMPare22rwURcki1eQ2F8JSq6xUS0OW7P++s2OXrRy9/X4ex8/pU4LgUij
vyqsHvwhl/gh+QzTiytNv2peqGj0YVPOKdcgQCfJRXZ5meM58Eix4NBj97QJxWKYqQik6mS0ueUv
20j6uAG47DqnP8PRpUB0v2fJnOwJ/Mr4QloNvZ33m1buO25NT8E9TZsgcaSfCAcMTsgU8fdcydBm
YnlvK+LCfPJHWa5PN7AL1PBNMC0bCG2/RQcZ+BU7k3QvYhTIb+sA+T7vx55hnEooNRoZTi1rH6wW
+398hD0TRU98hKcNzzZ90kn6Tu5wwpepef9VQnZGKtjZtbzYVjpYf9k/onQ9yzSY/IL/2/QfO/tl
Wmg6d31xq6RXztMlKbXYV3NLPRW+AZTVyJpWLY28HB6oVMT7MS+/cdYYdmP81lDzIp35her4FEo+
IgW73wUaenCIjiV4nRuAIL/Bk5kmHbFhuOLct0Rb4bwgkkhnauKcKvMeyhuKk9KDPWYI8hY6UXsW
PhXtJDy06CgKlFvQICPWZPKcnp0jnGnQa/eJOdl9WydkKJVoq61l0Lp8sQFfkwwy6FdgA4zsn0Jy
wfWvBOjjDL26BCZGR99QwIvwzdOkZWfClLWcBR51bW3qOmCZ9PRXFMX4Vjbg5M26j2NXYVSuM2DE
+Gs3X72Vjux3d55xp/h46d0roqq7GfSTxPbsCDGH3H8AqseVEz+OrCJipBevx/75yOEPnZGq3j1X
PYH6/b3SKbfprANfCpynT4Q82Hr7IKkZbBJAbXXzyhs3kzna+eeNCooK1WfGo8wZwQMzVQfl1apW
HxUA4YDkvoPZlTiKhk3DRDBw8+Bj4KmnlQ4uuG/2cEJn1lW+Jb1b1fNC/FK7qO4cTDRIrISQE0AQ
1wbaCcSowOwDjqQSt1EJDbPiKzRS7f8EmsPspTkMVE1jiBU/i5cKi5lFKxKeUt8Xzni4IrnwvQP4
osqdshIKzyKEkgw09lvkDcQaVPmrO/PBTCvQhLrX5aNiyi84Kv5jZiBHIvysSZnm6tUxp+mHUSxG
WVtucWyF2kQea7Dgl8STI7CsQ6j3vRYhbe2htUUAE6isMa1bi3xH0WfFEBIlmDUiI6+oGSrFDya9
Y80ilU5GaREctOfPCNqm5JC8K8VcPsgtZbcJ8y7oUeJz04+5a0LP18QbigPrX7MdptOTrndrxfBH
UfzCxlL+KH+R4O23dyHX6dKagI62mnX1whgv00PHLcJhiUWdT3jaIe0682vR0RWb7rIIFvcK9CYg
uoFKjVcnM0m2sW/tVylLP5sXpq9E7y2s+xuZOaLWyLk2tC5rt/wxLEItCkphTnFOcjLgJvWzcKw7
TEH/kzyFvTKw4c7Xrv0wYhqklMNMDBuVoA2/CdEpbNUpNfJ5M/bq7/R7LfigtuNVYEL0zOqFSd3l
FuSQZOXBLKRvB7kHQ+u7+7fci5/QECxt5sCLa0iv7SS5/6lNpv6L3PAGTiCpqNptXJ0Hk0hnfYEE
FIlaohVMK1sX8u31apbixkMCnXyKcYVkTatUTJjYzuPkjFiuCXNNPY0c5tTRmHtBgpP4+gP+Bxg6
rCZ0BrLF+2hBV9Nj2pagIe855+HvQRbxRO2e2E9u9MmIxMJykeFLWT3y7zxg/m1UKPwsbWwJ46mn
xWcKfb1U7HrRuQw2cYbKprZFPEtdoDdqI7t5sPFqSS/59UDrIaI4iJms6LWxHyBbnAXuYTFNipqC
QTdP8LKjQc1btD0mgPI9r4D8yIzhPqho28WGMwYP2OcTY67fvL3ld8ijAMSIyOzPsGlTSkqHne0M
4IVgVdmoYbdkUItyQaRODwcLOjOb+J9XPj+BasAZhPWFOINpbKmN7AGclAApD1gOOm+R7geGC8yz
/KkyaPiYePyBZ3SRxarMsL1KfDYgvb4QDtABw5nSTPX3FS4ByMzSRnb+oybSAnJr3dNE7kw+wHT6
p8NOwWR9UbEN9jmmRLiNA/MXTXm/BJiTYefQOtFc25bKbmgfvWnVTUffYfuIVWl2e51FNVmwsMTi
zcgiigKybR14WNt0qxynbrcPmqUnXGwaFTL2nFiC1ppyVzQtgIlyt2i6U/X/knZ7ZSvzlm4X0vUz
wm56XCOSXPhehk+FFv18tFu9qO2UcGHo7JaeB6/f+44WPNQABUOiUTEzjnDRKBGWgWDDsqrQdKI1
iU0ar4V2QEQlxONzmII1PGEGNSfwwsK2rKRWU+5FSK+8LO40k0GJNtgiGPjIFmv/4JL/V2DPzLN6
n5un2RBuoSK6RIqtjMTLmfzneHB0yMrCth9FeCYfwmjgqik4FMr7hSSWXnHtMbSrZj8G+afjb0WB
E3HBVq++NTep5B0L36j1qxymVZA3Zh3R4E3nCwr3AfFdckZ3iRpKn9n4WFEBbmOWDaOGilr5/JiE
q4eHydkSF0NJsL8KrhQXGgJlggMytNi6jGllG/jozSL3ToAKf0zxQmonJeVH8gO4ONFfW4nj8rJ7
Ju057QjaO6yP2lfnaxUBN68UJRVI7g0+zCdfSC/IZ0c623pz2XoZrRoK5cPRuZRYakkbygPSoEIl
MEwZ9tzA1vaYs552vkQYLG8xHqoiBLPN+Qd0QL5U0FQXtoo7swITmjqtC0/DOFb/7SDJZD5K3xP9
+HYwG+wNOkqe1qPqi387DIYWygAFURpZnQVqtZmYCesYpfwNMXzZZ+lnbHyZCavBbMY44t9eaMWP
PPEPTZUpkfQ7NTocsc178wnAcgTBoRjexL8va070tJf0//ehGhoFTFqVWM12HwMPKdd5fsiSowUJ
U76jqE7RFFJLBd8pyQ2uBOH3st7ERmacmIqOhwUcIwq9/XevL/BbB+KKlD8sPwmNwlH+82Dh32cK
c20SBREpc0NB8U2vw4YbjlaZ0/xhth7DzSr//Ks4qWVSvkh2k7vRdcIs7xSIf+KV6BOV/jYe+oqi
nUehhgytLa9iU9jCQdGhp1oE/DSR3a7tVnqf06a1B6atBvLyLOzZszgxKea6GOTMaJWm1bBXva8F
afxZFaViz+l8Gfdi6AlHLzWocRGZPvAI2sVeeQl7DUsKCX9Ay4XbCZTAy+K51ubseFBK5d5wuTP/
9KDVt+DpvfoHLAOWJD7UG/6LcvYM6E+E5Q4woSddN0hQ4+yW5+6Jmmd3afay+rHjpzxJfu2WUBwK
PiNfhC+gn/ARvZv5t+TfgjQO7LWEvbpJr9mTpZvDnbHss3jfTzjzY0g0T/zFe0+zPfaMErTSkfiG
q11T5uOdTasESBn3HP8DcuSwNVM/SzRs1Yzwp/HzugM6uJcwP2rWuJyIKemMyUxHoDcTqc9fta/D
Dc67oHOTulQwIfuozL9nCz20RsE3L/46Z5djLAHZlf/+tFGeXK0DRdg/f7M/94dmMgqZq3/OJoB0
TeqTT5mT2xCa1nZNV6JwcIUSUovRcJqKYi5cUg6PnGntoTn9fZEDSCsMQwvtAnHIx6JZfp9fXG9h
0cmTjaQNLthwIFXH4Qw8WCcbkKDv7yuL3b0DcnAJePbqLoIbheQWo7ouqCwg9LEZmQNvOPoPVy96
WxxB79y74JT6ie+wVOKagyXaIhCC7dtNhk+xxAMliDP8FlFb4gqK05VEijF16r/9pI/mm91BXpGs
gn7EEKS92V/f/InCHWrwXO9QS7lyW8uxcmeGokKmCipCUn3NKYEQsHpfdyz8N5qevxVhCosOTpvs
MICM2QlHoaH5x4wdcOl/pssr+bVPNghPBpIY/0cv50z+MvoOWdcgMA3GZQdkUehvRJdEui8RvzY1
epMMc1Qwo2NtLwwJ0IydcbWrqz2/dx2T/JFUS65xuvXs1qHgMmojZwhkZLj2eTjRrxYFe6Yrv5sG
+IvQhQRGUrIshmO4fO5kw18cbFA4a2pw23QPE6sDS5R7IValns6OGXw6nZjYucTE/BVlcrC4QD6r
VRwUIT9EmhjFokEdboMLcq1mCzLOQgozemVYnZjjXhr56Wz/BOKpsQlOtBcThOD1uo2HiDczmieW
GrQ2VstZtT16S24llP3u8JbYPV21ZVEyk2HN/ebIqkMC9vl3J3xGiXhLhMfgTne0F2AhHfsytM2L
9eOk2PpYrcg5dPi/F4UmIPocPwJy+l0dWcItSJ3wVh+46Gk29oDIRwjrX0qr0Ha/LkdQperBur9K
HlOAQ1ZglBgaFSTHCTPNZAVDiBgNLGCwF7ixCNN+MHchrxZW19xfMBVBqJ+a3LD8cf3X4LxcsFei
aiBkld9qInn8UVY+Bi2O8kWRcHtFfNAeNqaIBn3WqtJqGAYSwW5DvtrLDY3VAoq/xZK0IfoFnTIq
ZyKm5AQP9mY6rzt8d3yI2JbDSxsDUeUngLMi2Ae5vhaoCeM8QR903ebXW+wBer5czAFtJZW667/U
r9yC9veGwY0PUmCyphnfk7CcjApNp0xMUFzKR+Eu+5uCZ9unG65IeK6tkKSvGX5IxNER9SFoxmJ8
9A579GcvfUL6G3NIh1S2sP317/+So/R1in0q2JT91fQ2Ex4jCRVw9Mv+T4lz3dhiCUXJ3rsP7KA1
rIZC5Ujr3TO8bPMKz1TrvYRYHjZqfwZk5SsiHfrHykiVmQZdlK4WhpbJqjxJ3orD1SE/3PvHwa36
+c+uGAnaTW0KLHGpjDaSpSENRQYEnTIz8wUWH/vpLo6Hb2G71Ps5KIfQLIQ94Bc9gGd7IG//l/eW
RMjBYCF10b1JQnsiW6i0zkuGvIaqLCzqdbt0OZ6JgFk5TyGPO/ToA6qYkJUaPSG77bPd/axAMvcA
NCjU0ZWhjVJ1d8aV8P1UBsCSalE5jxXPasA52q2Fh3fBhEz85rOcmdS7m70XPa+EzFYXjlht2b3V
9cUVAz9aD5xDKzhUYMkubM5vthhcFRm6yRnILqQhtatQeNk3uR4BBfrF8gzWa3dxSiTMKfNCMWun
Ru+l/MWafRbh6ZYxMg0VBJuaYJM1ZxWDvuaLN690+GORhEpIiiDDOWC8XokhL77JMRWrO/5CAyBE
yvh0wlidCYuo4SqgPA1w3DhwALYu9lx5mWCG/k9QlEyizUFtEOnQNfcK4nY9D3b7msWReDVtO6Ct
McHtkdhCLuRf2/C/mkDmvrNc1Emib9hKP4OUcl4jW8iCU0e3NuhY7cMsuBaN5W1Z0mbzYdaFyDXM
kJU19rEXWx3CfgTfdp1rnwa4N/XOdiKVzllzIOojFD808xWLa/SFDnF6PLKT0cmShcBhM2tHmMoi
hTRF/W0YK6svKo3lYkHaLjvqakePcinHlqNzVK/KIo+68cq6/pUmoSL66v7Y2zYwLdfDq4p4AX3Q
qoVspPacx669p9qhF0QotjZHyjDo4zJstEMayQY52lk2bDud3hpWbxQA93l+xvtOyhrilaldf7Iw
dvFvjy5avXr0lzsAd0fzqZ2Wssx32nxSx8riRw30jooAJf1KLDWsUId0ChlR3yCri0cgnSlVya4M
AjBkr8b215eRCMZ5q84Umd5RNR41lh24xR3MQZr2D6BQAfIBAhRnRrtrC0vXvGQpWdxq9aAaJRpa
G5groLkckGmfZU0sIij1p+9ymccCuPMyfs3vaGAZ9RAZ2aUnLdTty/73f05o/milZ+rVnD8pX2OX
bnsapaCpVZLjicmSoCyRiWjWop9TFtR8s1g24DB4zabkWkHzue4VV8GiEQERHf7GmGlCDJodNits
BLP2JcfRwo6+MeffQVuFkQbq5k0qCYKAC3lSfi08CnI2dVvQpXiOABjfVKKKpOosZtGtmIsLhQpd
uD4NDM4eJVyopltZWy4Xmz4AeG81ig/yK6W3ivdWe80Q1SvrbXRrqRJa4fcNHVtY1Bm/79cYmvh9
H3qW4KFIaZ9SbPhYbHW1K5v9ciicSEVbPhiTNqdLJ3c447KVf4aL0kvvOxHymcIctTTYSKoUVV1/
tGHUyR26jjwoqNCO3ztK3lcX/ooxmcZ8kg9LlGTfO2VyZKT8lize0CNpniIb7XWdnzi0CG9czrfn
vmvK5zVOV20lPCKGsYs+b9y042dm0f/HknLiRqOqKSPcsLVO6WtFZp0i3O3BY953lTXniqh7wFoa
SvQhzEGhv9Lx/n4JjAdZBjGRohPT9B9BE3BefhAd2k0+rpYabHUfKMOPOfkh5ohQapXEaDLdPukK
NWqt/5I1hCxnxH/sC6vPJ2n8BRG3nZ3+bAPeDHwtcQ6iKr1c32/6z8X3OZy7nk1kt40dPQ0Awf/o
Mp0r0pCUFfmDSr1tNY4Dim0NDyaLdNhd8ji6NuItSegums/+BAHL8ggzuATbYISwtOXcV9gPkYxl
PYT57ZHFJ0P36Nv4weFJLaYFNNuKVT2bQcjjip81ptHQHAPJPC7HJE4CVQAzju82WLJBayx2jTKV
uhKFjrTkfGrHKa8Qs49ho91/z/BgaowexwVKaTO23C3ef3Da/H+2vgYjfO4cCKujGSJvzmQr3RFp
lJfiAbJuPV5HBVo/ntB7EItE5NYVFhTNW+kfM2T8G6YmzNFGhrsbDAKNaMmQ+3exdBKZj+Ju6Oo7
GYIeN4G2JJgrXo+Gh4HmNnaTglaze4ryUp3rY91CN9ubg/VR5z4VGWa7xPtsMaeH4PhH4VpLDZ46
X7NorShzjvGuSk3bJQJG3oyLgeGY2lDhhUS/jA9A2hgCFctzDGpI/m/vwPAQ/ya1IXzpZV/qqAcj
5U9qYrsddjUxfpO+6Boyn6SaW0jkstOsRpPzwbfkfA7DfHTJ4uO9H6GPCn1Ma4Ohi+B/+GmcfZzO
rksxfO3TSPiZVywS6IArEgZgsLKNCADlEIE45P4o8axApFiM1Q3bZQvsgoPl46asHAnnmupH2MPC
0fAH2nS29sZHneeA4PbkWxXdqUHtokN1kfZH5E+2PqhuqZkLJ6IBbVnvf6N950UaEPTkKop+aX58
vH4r7h8TdUOTvVv9g+5VvErPqQNEEq6LG1Xi0l0jZRY6302oLY/La260tYQvg96idju5JQcBbF3d
Uioll5hDXmYaIi6oZ/k+o/liRUHyBA9gaDP67UV4NIGg86AJXs30CdpOG4Yoe0zShaX9kZwEoh10
o5CPtygVss4qzfozfqnB3wYjQWke3TuIsBkmDXkG4BZY+LHvbBH9SrJdqODwQsGCsr/yK09O1JYC
4C62a3gELWbCCcvnTmBr/LoC8V+16qb1/VEvf1uV8wsgwTLR25hYprB1podCh546BtUyo5EuAI4W
zr2fK3DrKPpHQi7A7z5vzwxrXcs1B+WUYbYV2IGLBcG3vNQZyCjojTWdzMYjReAa8ZzeBozEtzZU
/0ZvFFxDGa62RX4Ua6uULXZP/KKQPjDhqdUdlSVdfXLKLYhaIw5B8xELaVZp+NBNR+noE+fD97n+
RLzR7FhYK0vsIr7H7MwKQPKAw3e+gA+U8PSVKSHFoyY2DgHZ4gT4WshZTxXB9nE4YeeA+Qh/sR8T
5IlD79i9cJnujqYUJeby8W3hI+plCk3ZGlVKBdld+pxs+8kH4cBtxjYcp1cwrQBaW9bM/iYrY7RD
FiLJFyMma8iXiBTUGNJx74/A6xMHk4/9JK6nKTGmkXtG6zTQZpu+7iaMg4vlV/k9ivp+E1i8tjNj
0r+1MSDUNQsu+xVc2DW2wAYPOL4WMUGOYs58MuK8KGWE1DRJTUXZlvusey+EMYHu8fElOGgOouj/
+JzXGmhN+HDLUXVibjYa2ZQzuQPVPy6KeJWzsLMVDA1BHTPeLW8mPGlcu13aU/lUae5RAYnt3iNH
29dJahn0ylknBa0Gx8mxsznPPK0C8z8sE7mdLTFAf6zyhMnSMZDgW8D4idk3+REmVeYlaKXqnQTh
Qt2Uoe1CGWjDEIfS9a3WGz7f5QSm9o2E2qZ2YcuLtD172+NlXlGwsqbs9aP1Mr7PZYPmlWqjuar8
/WW5BVRb6CFX6pb6bELDyny5ivlHI5pgYmzx4pYduc2Tpq/YqBLalI5tDcVJdl4RkXjejkbQBQ2z
0eFdKkg4Cp+xMwJz6NKpIjMUXhs6lRiOpVezRYQFWN+xIBz6xovJ1W4ERlu9ElLItPiZNvHrQETw
TbYTIp6csUK0dvU0fK9wg4/J81G4nYlVpPpMtfjR48ftN10D9n0heXBN165nRomuXGQJLpuZAeYb
aLA3ng82M+xZHpeEofT5hJ8PWsvtKhI5VQN6j8e+icv2q69oequzZbajM3MyYV4U8xBxTw24XDAk
5bbHnHSO68AhuSjcD/xowJ46SfxF/o2/r3zM8qeeiWV2Hn0MIuSl9jhTGgt78rgqZPZ1ViwB8YsP
Ld6devVm56MtyG6vggPVaBp6ZjBsvufo3hAKslzuecTatBtOFG66EJTdx6s819rcmMYNL4Nvq7je
kKg6qd4f67u1FrC5Lgt08w7b1vzixd2C+PevJL4NnhOn8t+WPV2j1t8Qf26kOTN9inqviqPy9DbQ
QqetUAJpTI1sbpa56qgK5N9VAzJg9PmrZE2+RH4vm86Zutg6l7Q0vAKTURhs24v8hQcADdKHMbUg
O7JtrfYP7ie/WrFLG+XpO2Pv4dA8LsBdhk8DEPLpIwas5KYOikeS0BccoUdJlOAek45Bky6j7ViE
DM2R6XTFZiDniSqepqCdFDI1zKsJu22X9gHzqSYWtEdmF3x1I2pwCRcVPbslHEf/G0V2qJE9Va+T
n/9gDzHTz57KkD5sgPuwKEh6KTC80mRoMRoOIwpH/64M3fuW79oZlUwYx6VqTlgezEYo9/jPXSC7
arjQyjS5t/3hXSjqreaTUrb4b6XDwbR610eg31m+ykS7vxdxTDLybVXZOex7hRJ7Ztao0ucfy3Sv
wSbIM9udXsthavZwaDtANZZm4j1AHzB/6zeZvGHPHjN01mfD3HuiGiE8OYH30t1VbufexhXy0hoP
+9MCq2svCad2itRKnaiSCNUmtcweD5erGq5Uv89Q3qIuvisZL712sOh8t01dvsx4lBh3dceareR6
N+iTfFQrYYWukg9zeDWwPCxq10GZmbuORjNPK7M0lm2DsXNYdpb9cEOUAuy81E6XNMMhta/jdpWW
66Gr/Ss1bp6DNhQJaniFw0XZgm6dD12EydfpHYFMpcf0dnzB/3bV7CGI/JtqkY3AkCzCEuI7ph48
Nhk87GL1Vhh7MXK/Y2H4ONl61qepwTlh2M45my1IJNkGQymphl2qR82WcMBt2vL32z4JVG9bvTA5
HcAWDL8QrexJhwpT8dE1fyDeih3HAS/X3DHNu0+By0hU+syxJWpGQQixk/zzSbDEZ/+k/WjKhOim
fOk+WDwFV9FffKo+KhyleLuvFMNZa+umAClsQkAUjxq1Q4RSodKiGTsXOv50akzfqHi94jjI41Mz
/pKYjdrVvVzDqyXY2ak3dME+AEHfoxfrC1yBoMqp3s/WldW8LYfOFI928OpGqoLNp8wVuXUWGvnf
IMLpaXnUOuLHGUpS0Wrha+d0UpGiqXrQQWUk9iuqG+SMzFJLzqASO6h59/TmGNhD69FvTGLImWSc
Q6oqQF1XnJ4nv+GsclD1C0rvqGFJDrmd+3g7ys/30oV9M5gGAISOknp1NyBT2TpD64T0dyQjNb6F
Cd4Ev8qWXFApDOvNPWXyBhze0c7K3ygo8n+qbxSVArpVvUJwE57ZLc1/J+5svXvJmqJvm+TF612X
l2bed7xLHbsCz/doV/yG1vRL+qbnAV2gb42nXYX2y9yToO8kNsZIxE85c7lUumOiOcJsoZ6BfwH0
3bVZ75BKjVdbVRT2EbP55ManReSz0IwUX2WfuQaPFYzn/BrsgiLxnQOeAJwZOD/hEmGFWfmhXi3K
MZGA02LmxsIZMIxVCaTDZcbTzTELFsGSN47PzC80FSLet6cnko9Cl4Et4NjCU9niIUbgq658D4Cg
5EiBcbzVUkWLV2/gyMjfA9M0FppCt3VlZ28V2CjkOhkwBJkMvCBbr2n1wF23LeK8FV2OMKSKkrpC
Xz4TNQFnA+80zmAVOB6un/nwCiUEShZzdjWeqpukGvnMcU1Q2BN+yojV+XwT/+USAHVLvaEgRZ0m
sPmvQgPnhqKFTG+M75jwKGF1Vk9TJnAgsEdyrl4FSh+IonzvspXg20mXz2QsBCKlxgw+5hFSz8W7
f72nHkHQihcJ23ZtGcpdgvoRxL7O6YX8aJqdBUSi9FJGVSf6vKfZrysg497LQIsWUS/HcxYe7cC2
qvSSvy83XZKy9BbS57IdCvnCkqbFjcqxBgT54uWjYq2K5RHgZlJDuLmRM33jinK/dYGkfvvIgXU6
0uSwAtEtToVA5H+HoRnF+ssTfijuAUkbwQjdZR2SlIEjkqiHZR4Vw9A2oo6Q8DA7e59Dj68iU16X
4sFdx+4FJfRuXVwxlsqBjMxqJanIAtZbV9ZMWxdY9x2cwuCJYqcYCcY/ZiCwcMRa0BYBjJvN43cV
WMwSfECWkuLMUrhBEsTbBaotKzBzRmZ+zmDTmbEQ5c+EckMxdZPL17zVSM5UdZR9LA2Ep+uOtpzd
LYqZIHPUF6XTK/zMS5d/93t/S5DXO8ZNAJBuPq+BKVivfl/H6kqI4nHMYQBYd4BO3182lB2+pO0b
rGP/f2sfUmgwuG9Nf1i2TctYGgMzuS3WLk3IFzYlzltbrI7ZIr0uxUxEknQVbgShy+jw3Oqwnyb3
MvGp/TFLbwwHjmPWRMn0fu2YGMAYq86rM6ENUenop+MtKmRCYVqsS4XfD0FP7z6GNb/H+7JZE57N
lqUv9k4Pr+i/SayZPUmNhNPQUXUhumcLutXZUuRtekuRgjwb0tlx2lSmJ4qZw8GB1alrqBxD0NVM
BK0SGSZuw8fl1R7VTYBN0aGWv/f5B9yNrRhT1ilv4OweS79LOvYGJwQo910cx0eyplnko953ZzFX
722l/KmUgmbBgjn5W/U63TX4MWaA8jDQD2QuH9Z6+Y1nYiiJ41HYEABYEmzP5tCe6Rf0QkJSNbZF
IOPpFJJISuIXCXtKYuO2s0J6F1TY0T3mDOWTCf29dI3+JlljuuzXTBoaOFhwMP86nkRJukz33OK6
hlPB9pVPLv9g0wUkzF/jiAcITFlVJ8isTXfuy1KiAvIXF+1YDv95MVOa1Z5GJkfDQpl8HhQZ238Y
Vpwpbhwy+++nZDYa3xj0bBpXkFRT7VZyTe5qG9jUp/Rkstum2+LHqgz/5iF9UaufwvsusGb5cSWK
Jjs/EVt5bulEVB2jI3u4oTRc/Jtoy2EthtHFvQ1gHDPLAk/kvXkT9uCrP0wtwMbu1TjPixOcHLWE
0ybF4d5wzz6pAdjBssVvpKPdK9jM5QWzU+MgTBdSkRW8aOqvJz1LrrTsz/xblnhu1hQGhaalplpd
pB+fERLJFOlB76T3lAmtdFcr2/Ng/7jIYbFwUv1wGamdazrkpGpoTJaaAIfLUZq245dLwpmNNEKD
nCQPahZ6stVirbMsdG6m/GQL1I1FZcP1pMLPj+IXJMaMrOFdhPmB8KemE7l+Yuqq8Ke3XRvUJkbQ
XmUMtws6sV9ZaNswzimLR39L9T4ApL3XMJbrgOhra5yj9jnCKJO23BugSBmq2UQo1W/fvjCHSMe6
vGzLN+eRPUUjtOFnVNx8KPzD3pez9youoPqEMguPKSmUCewd+1PZADqRl8gSDeNfUJ/NlicQVRfi
yMHXgHGF73UvBnCKm2NsZHdXNkmDqXPOVHjaq2ZI92+57I6Qur0FzFCC7kDs6EF9ijHctNXLDS7A
5pjnq3KOtPPFjIV+34vf4RZ/Ma6tq1RUWQJIIARZhPdNk/X+xd0raKQKUQIsl/umUcUYMUwKR+wv
6c71+ICGKOTDL1tczZDmP79oUa9SxZbUxTJ+LBuYaZyV7qjPII9cVrQIXISwDSbmAJEGcYqVSDhc
0nohG8hvjj76T2IbBhnK5isI+2gQaQrV8mYJMW0uH9FR6TSG/VbFZYFxyskaLPb9qj58mkLg0QEl
TLms/D3Nv608Puc/ROwVq2KgtxJZW4V2yZ7DGcY2eVG2GBNfjT1tW+9Ai6kJIHpj9SpxTvfVckul
hmeEWOwL6Q9hey//l6uGKCbkpMSM3uqNElZVwRtEYKhZsOyPwgkoQl67jCFs6ls4ttjvppexJGd+
tf5bZ9tsIN4Gb/lOcKoeF2Qgmlu0aerPq9xdKun/mI1g0jhkJy5uLYqPLXSMBpP3xrnVkxFnpDpb
kVRrtyzNLg8QBqzHo6lNEWieGujttecMiPBZ80KFrC+E4uuitcJzqEkALosYIe4FysKUX14tsP1v
BEDfeAjO0CTuBTGfxApxiSBvbem/5urJvcZQG+ARtS9YvFHJXdRPFFGYUYTnmRbtnb7mvtnr2haJ
VpNLxsA6pjnYFjWGaUmd8KTvlzUamtEPlJi9bFfKaO3P68+9m2NekpcCI9CzxgKqlgOrtJZ60X3x
28qlZlOeUHfnVdMLxQ1TEBE8n12J/XvgkWW8hFJNbwKRnPchOVslMMr8uBbijWByS7JGrs6JuWR4
XRWS0qIHmCaaouDs0OynZ/n1mbrBqm+SVUDEPdAHzxIx7EVWWSnkLfuqN/aU8ORK/fUTYo8jRhAU
XS+I5L36aQGPCCHzltQtsAftNm/Q77/LN/tOn7CPJzEMclf+136qsIGK0V06NVxxInclIUtiRNxl
Uxm69sUydc6CBpFnIpWGsB4hcKcqBoZ9y496dZYE5HNqnrYYuB5QNh+9A+hyeEVFP0JGbNnb0nuw
XOpvgI4rj7UGI/fLRFdUA7D2Q3E4k+N8D1V2hTsiveJwVqsyUVNk5iN6KXiCgUmtqOuxXFk5ic4k
zvx1ADYp/ZcSLnWPOwqtS5jgKyBZ93luKUHrOUaZsWw/dmuu34WNAhpoi+IdQuBMm6CP1Im06eRT
Rw1u848R0w6y5lARaY/S4XPf2u1W6ofmAGbuTMM9dqSn+2QHajDq5zQfcBKCNMPAFFO85akwJgXE
lThp2K89RJWkVZFIcPkPCbBDliERMLOw6iNeDKp6334zoHkn9qirqhS1vEUT5oLBfDazOPn6frU3
xwtQkI5N9GDCQax43O9N+YuctP8nKm2kd7fG6TLe9j+RyhSHJTaWpic+nva3+JsRyjQeA82JhUE/
y1PeVbVvf4g0qcT7CKqixjWYrcWTYfb8h8niHz3MGkqc5bYmKedHD69Pjok2Omhosjc6zONvLNUu
GnPq+zuvjE43vJrtsqOPIH4Lx/aRehIdieMb5dixNlr6HfeFuboN7qwhZ7EudFGs/4i5a9mjXrkZ
2bkK+NNib6c8X69KeZyvBMISEYgR5xPnM+0y7yWi/TBvOm/irewam+IWbia/I6WoPFCkORzYV5OA
MrUvxbsptB3umqQErMrrkwqeAidKWlKwPCovxoajBdH96KRoTrSDuy10nYOOdW7N7ud+CYFRU1Ai
UPUm9/gQPm/8g/uCNp9heyIuJbSQYBeaJZR/dTqCkOoxaaZQXm4+PcL8qObD9a6i8PlJjEAJWzVs
TGnDxBXIsXZr1JBUwXsp0Mj6EarKGudR5rL8NoaRa/IYyInaG/D6u1gjioMnsT9ltrfEGO1E9Wqi
2UP1enLcy8xVHNRsXP3UJNfMw5x3AAXNOuK7lmPa7ODzuOF9ec44+53TaKSCwOhmMEX4ZgLb44eU
FsRJYAaqeR/6pwx12C3XFVKusrE+DaTKuNQK4qNH5cHmSY7l6FphyxX421ktlJP6HuincUabY5Xs
bHaXGnOhTKBtTuJQiZvSWLIFh7OTqvLV5yc1J0zZLWtvgEy6ZQGbwjQoXskM96BQHpLNYhMXzvdw
EsJWW3T3gkyNaalJO9Ch8kVyQkbglRaezh9fWfLdn/vizSQpNTr/1pIzicc91yU33LechEMwT2iM
rWmFT9mBxgqGu1R3mHmxDBYRX8RSXm+caa3+cXlr6k0lTjAzv4ERbOtKE1E9yHTsw3lLB6Y63rrE
Ck9iF2f8kwM4eCnSS+aXg5L/P+hoslTvwAXIXjTmbakaYnkoSIyNLgyS6YNDJNeKebHQKa8LZEKA
5kC/u5IfshsWKGvtB+jR5WkC/PUJSVfE2tfavW13C7+NshNoJzip3HLMR0hofOOxddK0d93DaNeE
Yp2iyxEA1e92vzKapi+REWHCCVUHr/P75HahXtPqKKPOxvEy8gIj36PP9bNdOFOYkkxOjQY+hY54
UY86jUta1XjCOw/mZgHlRjNkvqv0ZwJ0bN4l8S+2OkxmZufCrivGvBqbuaqhlh7QSkAp4xgJa4D2
QLihbICpOrWTpIPFl72tLXPqViBR6h0Akzmli07mUcl7uhwmIdSu6IxmMQA2n8tSBJ5tafItXGeX
5bYo7FtL3zhitpYxIyHj3UIHG5m/jThri6pDrv5mZ40Xya8QXu/kt4CUuDeXcKRdcRNZ/2gs0YMZ
8CVWMsjGzfdknqq2AtWogQ599rVc8OXgmq1OXpkqG4ZSah06d4CQoTgtiIRcVpfIEFyErsR08ioy
P4G01ZBYVc0RcZ73rRdx5rqk74hfsAG8OQGXTDj8/jftiucZUG+R1DAbmNsmNYVHCijR+hFWbDZn
zfY0nlnOD+nzcqRKsuc4379fcHsM2NW1byqK7Twj7JF4w6YOdIkvz7mRNvot91WCmgFUoeHC4De6
dFpiiNWpdlwJyO2P2HRQmDP3TIQEUeoK/OF7hJ11ArBFMfBT/SbBTNSNWzWGS9o7w+zw51Gf7uT7
UaCEnblSwoCvnNTP3IoeiWpNDsO01JiUkfQPAedvDpz89MPd+gVXWhV3lW7dbUher0Knk/7ThVrd
ZUNC3otZXsZivW8rkkzMOhW0evpKzzBXzaKRpvLrSGRt5gBL35sY8R7du/7E8nC4NW5PVVvO5dM7
+k9AU6bLjzJszLPw4we8cpJAypLy4/8TOuNRtnZvk6QzP8x404Bq+r2orXE2KfBno61nouL73Z9r
yUDel526PI6AdVXKYi48lqZ+OxiONskCg87JEfhyqbcy5GURCEwhhir+Hsm3a7zJ3gdpgV69w/W6
v5fQsT+KcCtsO0AYdFQeKb6FFTnnZcPl1TH9WKYDY8OSUTb3v6BhssxuoQOMiwbkgrJ7YLIphUzJ
AH/bSyVKnvzokQBvYcHFc53l5fUwGrsp8eZyVWA7JpWQ+8C760cHgRNWKa7lSLxvvi29q79Y6jhP
AybPxJ+pS2UX/2a4rHqk5B9Aqtd7sS9VP0LJdfl7NkrxHAEn53cozYgFIH4Rxb5dCsb5pBlUrrm2
MAg3zt3S4kEknGi+WG74XcJpEWgMhpIC4gNXFXDBvp4WPplUr3WQABEHiEs9nplLjdSHXsrxjuqf
cYuoikFI3jxlaqae7ift4hV1uXug9LeBeyXpwOXm7ehBzAVaKMBh7RDvnZ3oKgDkSCEGuztyScW9
22KQQG2TeMi+hHfQ8CXNL/NuSv/rO19FfN2yCbGYzdu13vAxBUFjJObq+HnpR1Sube9krFH0Q9HS
Com9QfARayftXTz6trYCLvUTTWA7myXDIPOcHEW190dNj5B6P2UBcX5/2tuJMhuKsEyZtbKuc1dm
L2nNcF/0/jsY17MK1fhc/t6Q/VmNaVLZuoxa77HMPH3/Vebgsiz3//WryaeL3byvyh5UZh0qwwRo
UBNwAMG9lbbrmYRost9Wi2M7amtEJzyJkLda6+Qc5IeJGcN0GtCsdSSdAP9iZLCctnVciTwg4j3u
q0yggPpB/GnRx/LGiL3otRVWCZrYNwymWMQ6+scaZYEjnsmIFlXVHIpDw9RG88wDq9peSTpVBKE3
GGYS9511UV36aQQLTS+3eUUH6pH/EYHvFgVq+RFac7gDE1QXfjNMIKd94M8S5eTP2oNl7xxOC1pM
sArPOZ7yE+v+jVgrgyvvEztnKF9VL1Qpu8p18Jwr7q2jIowlt5/fpTiJAvpuMZboMMWoNEbVhKww
YA89wwGs2pZ2DDqb0RGvc8RBgEWE6N3U81n3Aac6mQ+Has5BTCL0lZYwe5hSrAupJMkdOBIKZFWL
OibX97cU6yYIh13JkHWewZ6Vr03S1VKjHxqdxrwWL+W5kvRzwZYsbm6z7GJApEVJF/KnxOKgJ9pl
aS8xinqgBO2JmJjLu9A727uAI94G5SJPzC306R3pTcybZXUBwXu15kiIfR+8JoYFE6klHW00Dv1d
57Sf8zvmpLUnnmrqWzYsk/kUwLH3Ot+tknit4aLreGiCJ4RIv92Pap6n+F35iCSPElGnuuGGv/p5
qgSWFhPqeHM2I0c8bnmT7yBPJbutwyRHZPR3T5VRcLKMKMgq4cZzsXltyTfI8CKHJEaLQWHSiYeZ
esZv/s9fLk1S1qLFaEWdNKcs0uirSJ+rkzG9NVkrUu6S1abu/yB/k8ISTCaNJ6MePTeWjvD6xbNo
wjfMa/RogISNrm8P27RHJXtkMsuxp/LyKdTud/AjOoL/PEu0Rlomepoa1e7KO2ns3WFwHFih5bN5
UPAaaaWcm8VR4/mdeQPeRlcJVV8SOjUutcYy/KZJcZgEjzEumpLHyJNwtVQ4Tkk2WDXM9TXRWEFv
8TGrH60vYvPvV65LOy9IM0hJyO8OZ5n1t8z7rEFb9mkUvBuiN/drSpxBwlUsSYXhmUSxwhU5a5Pe
hKf4Grkpsm05a6q3CiDvlVWB4FQDPqtq+PjYRvKiwIQoK6Xz8GfDujRwziCNBJKSdYQqODFTQhbm
RIimopCvHZYONCLWfH95mPDHcosPA4yi0HWo6krU8oEdPjltEP+QRlVyj2AwRVLhhBR0nioMdUdl
fvDZK5s/vyutgo3ufM8trTKPvY6JZSGtNvk6SAMNZIWIU2S5pZNb7RSyDtwMJZ4GWI3SNshONTrt
MTe3lo3QGvw6Y8yFUw2Z2kyOGqmdUQZtsQ0GhAiRRECsHv+k7bQ/yGU4Ta981vyY8fvWSCGqeF5x
huRWSjx/c8v2pHzoQVt5yP2PXZdJJ1JtQ89lIARq4cp5sA3svD5wQ02t3JIITb1HHhhTYCKrThld
ETDc0wXUO67c6UTXwXVhkUEHbrfrYWj4NpWDRTu56qM5nbV+peHWf0sRvd7xsKfwvLa2H+fkoJMw
0hom83LR+vzWjnPUUajECMO0uq1R2OpWmtPpnU95A9Ea8Tg9a8EoIk1RL9rMI4mjTrDy56FNfZ51
xFkeRgyfVhbMnVBdl7xeoWft/o+rnaEyXUiPnxlDsUCl9oOCBvfX+2MBPd1g6+TB+T9/mMpSL5ie
913ua2FXtbI5HgzWCG2KHLLIbXk+q1TGbmw7IjfJxnPAuLkZfaBYYMfTkVzXCZkJoQjfz4wBLOY3
oqTk6EhK/OSBg/ekXU50YvOsEE/pA94nUmvja2kUYg+ykMciyDcpncXp7tMRgleJMRn9vDsI5zXl
edzHK08hOCbOT4+Eqt2E4yiMh4xhLIr2DmRSX6DW799gXyIrrc5JgmKlQ6aBj6Lp7DtRKa7U6jKd
kSQ3r04dBvZDXzEaz90pCP1Yag4PP++SbHNLhHFAy8uKC8iWqghVu3TcPsyjJz//qTesiJq1TD/W
w6Y3Tgoz+g+9QkwbmxKiNA4pC9uXqfA3OpNn0MCIjEN45goxZ3K4kQ2p0xXuk+Q5czXld/+wUxNr
WrWsM1CRPun+HvRkO/mGy5W/fIBDAlDP6ReZz2kGygr6iXY6nuzJgoth2DvoJD6sMczwmsYm+PTe
+cUiBjOjLipRei7RvPVGXUPdav+mPIG4QSCV8peqcEa4aj3RlMT0tymlcotWooS1mb6Cel4JAO5k
e2mhHCxg1EwnHMXzVydpSHbFpx52QQeIh204IXore8Ncu8OHP5/l3QQzXvx1e2k8KyVRx5SBflZe
ZqzD/O688OHF2OXpScy8QAgia7pEWb3ho15iNUfbq9gh3HiTSzAE4verJamjH+etAK3HyNllb8eG
UcEU8al7Dg+CICcRmuPkneemVEE2BDkEo1TgZbU3MIDJ1XzBJRSMsjdl3O8gH6ATrpRwVUjKyis2
XL9Kxr66bCTQQL3ZRyJIZfCcHQIIB9Ok3WmpHR9wQC0/24Cgw+tAXneeak+gNPrZ8uDvJE7vCd7m
PrguPxxoxI5KwrP18j0QnU13ye0ujHUAq8j06fw//I00+qUnwFFRV9x4QgYnhP2DV+lpURFxBkJp
9bGKblFuzkjpXhatjPmf4sTaM4nlhDhJCoo2lzd0NLNmDa0zL4baRoMtYmkbOUsgmRnonk9fHtrp
Jnc4Aka6nlo/0/MHgBH6+MUD9EoG0hDQYfSvQOJ88gmyf40aIGAzbMNzKFqNQfGNUX+ItLJhKROY
JaqafxJxlhQX0KsblrIlFkm2160usX8+4q4chMsbpHL1daYwcCAd4bBNrIYb04ZP75yjXa3YTs/e
Kes07jGHGNaoQtvy4322B03Wg9VBY2NLtPSe0OomJ9RNDEoj80gRf2+13Ux0lvANnApHrfuvgGvg
TdJsJvu5ItBMKpDWd4dib9cVCTk4xTbUHBmBjHwbIFv8cDyYMBXH5ksQdiP0weBFC1KJmaHP1JXr
SqErLujHwjsGa4PZ99Mx3PlyEEAyFaOLcPOmqaZw45djYk9NcpdASx9KFlMRG2fLRPDOaxcDDnkX
nv2XejXjFWiOn2TWUYBt6Dw/COd+m7QOulP8MTRMVP4xo37+cTsVQ0V8/2FR80lXls8Cv/3sBInj
sioAt6WDINgHYCBK09kyWCL9t9hyDizZYbTd/prGK2PZJdk4G1IetrmpkHC9mW0V5XkcKNCp6dEt
2mjPz2k/ZhI8pZQDjAWJ6eJaDAgxjPsoSU8knmd2HCH1FPqjEO2olzN7PJ3UxDih7h60nu1TUF5S
MQs/Wp87SNKHSeb0aZdIQOqWIxEOJcvJdRZZOXv7mglNOyuvNVCLjJVYqOZiwKvmOz9FSCwUcSY1
9MXlawkgDjH6x1fdGjK0lnbVJidZRDizU2iy+L2La+XbRZ9draD+5+iW41dCozTK8r8NWg9HH2Mf
ZWgAhHo+If/O2EwBXEV1DFeiTGSSZXXtoLzyQ3pjxyhyflM3PIknSjo0oyCbno1ctRB1ugbzeyW/
G73P6Id2J3vXGMDiWgplH/iGwU7DR7b/aTWDMiL94GriSrTvhd7QKhbynwGd6gUcyamA5DFwbtRt
1Avl/tMMvM7CsSHgLkn05d2kw2WxcU8z1yvZzotgGykd0jDoXqwPDdAxd6tmuZcD9EduiR3i+bBT
gYED1YezQUUWihvYB03E0zBkYsW8gc1mF5YuFIYZSm38oG+4oCFDR+QoxbLqMYFF8oCrjlcwBeWk
HGp2aBwxpcNcIDu1jLALhjHc868NwZCjePUTRjMn+F5JXdWIkfdpBnK9W0+sHd4a1Z2qCL/xIld5
HpzQPxZOpv2CYni8IKPiPXNehH5ia9lrgB9XjMu4dfk66/QwzorDqKn26NFSqAWW0TRSLiHI+A7F
+hW/JJbCaVwMrXJK/YoW/kWFz46H1Zon72ipnZC1iqe0AWPzTn2Jqc1eHHU07zYXYBmwqCv4zJC7
TNmJOguaTscrhUXmm/zCqGi7ZdlcC1bzN2TJSRRZavJrAU8x1DqHpppKvnPICw1efgMMNdP3dzKE
6oa9u5sDIALQUSJFKlAIEz3c7IVNp2g/pyb9mhAkjbgM7sk++60j9aFuSKeDFlZR9nNjUze8wlqZ
I1MeSBYZMb5yhgR2lmfgnVFnj/uzovB1T/J2Q2Un/vGkPoMf3WX3UyK02bg+ESTatT/llwANHu1r
hNHhPga12g1Aqw3RGof8hogZanLvW+4ltbKgqhpEPOm+SyxneIFpJFOuvQHtccGWUB0ndSwFKXSk
23ldemo8sNHyIlCTw0udLxUuqbb2vrH8cr551Z6mh+HGPFNv46+3AqY01Jm/iCnudvNupf6VCauv
GfCeaShFjI7E5Zy06QGOsxGYgbHoa1kgchpGsScZurXFby67A3sHe7/F6Q8ukbLXCbngaPoG4luo
Eu1v44kk6ChMM0zxz98m8fNrPQW3CwBfhITnBF2cCIJ6ueEWKi40zU+prM97pyZTyR/4K3066Cnm
UlCSGvJ5m/APgmU064xg4EqX3Fguyz1p7f+bjasUo8ELbadnHOQAm2WWtKgz5zu+2XoPYpDbJHka
OwfGrmkn6zWpwqxuTFqtSWLtLEODVLq5tMJpsSOyMQL0kjMULVCZQKdI/qMp/91W5os4bCw9U3cG
TRyXa/G4sDfXjrPTAB5Gi7ZfS7q0hEs0nAmvoa0o179iYeE70R044GDSoJRywCBSx9b8oIn+B9gE
52jeJ+ZlXKATmOpL7QSCOK/M6gWd0gBSR5fcVDxLg8/6eaufolkOxsI1uEmJx8vGeb+6bCa7ID2f
FmXNnxJHv0e5K+DZVsSgDnMrIGHbmihV6PQry8WGw80LnElcqr4FnkYehtzNeoQCorI5GOdwJTwV
CYvl2QZq61bIELTGabjCMI5M6Q1JaKkDugoiYlhik/e7z7pnt5kdbWZrD1BSfoEefRF9fjF5GQdK
MchM5+n2MrfnExNA55jVKTICG7JytM8W0q4ATxEj3dbtdhoD5vx8cLZjbmFXTHgVhpE2zD73W/sw
LzXKiMOyFRdgHim2Z/6Rdz+RxDj/CT4jTCb/mr/xI0gP00Xb46OdZvo0NNgmTdSs1hnNvUt/j2rD
WJtrCZGEGsbJdWUQNqCWNUC0Es0u0QfaakwmBVdP5xair7DRosnoO5kkqKBg7NKrxV5VhSFgwrmF
yAM5sdIlMvbsR3IqsrijzsIXL5oXhk7cJhvSbMTlgTVkRlfR9b1tuJ3dBUOyyhRLqp4aTq2vvXg/
Yyjb2rJDOcoRFWOlRIU5tAa06uB2VxYQ31ZsozyHS1bse+ar5mrDh9SabyIioXcGJQLNITWea7Ql
YFBEOXRDxuhnZRbIlUzDBIp7verERTOFBbJqNUeaI7VK41b/SwA5b60XiNpCCv0uhnSDkbeHxIRk
N1VMwulW6/NZ8SJcnzVcCDqoNxcqstMbLoMW3g4GlAzzhELesznx2JuALZ5s66V4UvnGl0I8pO31
qNmRp23LFozXCOUqpAnAcsK4oUwbgjq8VoddW2ipW+IFNgCOk7rQ/x4he2uuueMQF8zDqcCdDB61
SI6J8Z3Sm7dITlkCUA1GZWV022eiV2Hp7oVUHW2Vo6EXb+Y3EozbvpesYdYwC0zZ+zVuZ2PhFLjz
CPWf+v72R68zTcUythtfhUQfnPZk/aUS6Jk25el+VWyj+jXOB5ACNZrj5sZlkHdSU0wbSn1ABdhV
GPYjUl/DcPHELxpoy+xzPDDHoPO9ZkAnpcZPIX0rqZrDAn0Ynhsjuj1nYvfhFwm00of4yrvOeB7s
oDRM0o90Lj3XWbvDt/EbA3DsRG6+ci/kpIgeYzt99pS20A5PGPEwyhVFZh6lZ1VdzVfyBXHVIeCD
Zc3FJ8K3DwxH4XgyehXQnaPitviNKUHo4E89IlmWzSqVZFO61a8v/GNM5VVzJWdXRuBh8+P5ExaP
G1b7LPkhOLZDeuRii1zdv0BkyMboG9NbUmbe0pl8piKMdFdkUYmXVlkOcjwqrB+V2uX6J1CAVliH
iLcdrUqd5bu/DrJr+hJu+8igutOz/6kB8wLaz8BRJ4hFwhvP/ah4ZGVzbwspDgJh65kgZCjx+BFI
PzwdeDVPXUJ2kaOD252iq6ViDOHC5IRVzxPHDxEBSF0QvJTEJyFr4jUe2CHc968BKWxOTZXBOGFO
0EGXABDQ7FMb9N6SZPrO0IVvyJPTsCJ1jfoo1fnh0O0LDkPTQtKiViEyKgWoc+lwswh6EI/H3+YH
+cAT54ejoNaMVgkwTO3WVwrnzqmXFTtvr4UaxDUACTfPYe1rH7xwu6JZ9BQ7j8GcHnovIRxCZ48q
GNL2alKHuznxBBlj08fby2ZQ28iLcTzwe7GM5OoJDBmeZAy/aWcx4DEvcO9v6AhmDCJULc5BmjyM
YWG1uB5B2LysT9O+FAzcSR3rpNXYNIH61uaDCYIBhURqd47XGSRKIQcl/xXxnzHVScippVE4KYzh
VPTuzzKOWs2nM4T6Pa6OeodXIdLfo9V55trtQPElCvQsQkHRIbm2GAbhfYVWdohapOv75ROf7Jv3
D+J3b/f1+Dyk2CkjY6Oa2T72nyTpd01Bngm81OiGsae29apUZliMxkLsBp1u40uwRLtQBdZPxMmW
WFjixCZATmAc2CTwAHplcuistSwh6hNdvT3XeLJZmrdJmbog+37mf1YdAS2srrfs4tZI0jlNARLI
XTAEMpgxtcYir3G/JmbowdvpH0bHpc8nTHYj7JqIqr/ixxFr0yEBSNHIb6+Ryzi4F1JlG7yhU3+q
cmXaE01xcF1j3FbY2Lx7qm4ugtb3IHWYxlT9CMjaZIVzyDGLSu2wLwRLq3jg0CqV+PfsM8wbpv8u
C7uioWv3U9Cs1IEYP2B/sL3lmpBS5UoIYgfXDWkTt5AZO1ufdz+W9b4K0ZhWIrYx8ha/rvdITd6T
x5UC01qiEnuH4Xo2b02dZyGvJeRN96+DnG+Igth+HINNzYTPGkwrPImm1ogORL7r4QTXG6iWkBQG
V5zS31acXBGY1ZIIZkL5nT8Ymo3yY3LuNtVWVFLVt29Tsyr8dMy+wv5ilBeXSINkci3N8tYIY9wV
Pn955FvqvgvIiuuFuyFpGfqtffyZ2nevsVpjeBmVN1TEn2BEQZOPIXlOd9OUGSNCbJ/+srRwYiZf
qU+c/DHkNSqK3Jk0Mb9JDsfZXKkd3JBeaAMnTJmx+pqdWIUcASk2Rrn7glCAhb8BNQOSfnGLuLz1
K5MPQ8u4R/uPwfGrBJE+6qJhhfhcSDvMNYAjfESDLSk5ObP+YtubLGRUFIynN+IdiI+4Z1Pw4oaH
lymjxMsAorRx8JX+eEQIMiN8vCBd2oFYkDky1vNZXqHwHJf/KXZ5X9R5N+1YvsRk4akuBFWENv/T
1Tf+tbUaWVJhIVXbGgaI0VchldsMiQiUVKm0V0PP7uyrWcWw0pXxMHF9oG7R7SxEhlvhPhsdaT/P
/26SbEoxNROnb7QnRdtzHfXdfhK5I8xzYqVC7lOkvSMyIojYtBXlZoDTIblKMZSEriB3SPAu0bPK
1W5gz17ohKrh811E2c+QyBTvPIZVViHVhVAerVPe5eGttbyVjbwGmt1wniVb9p9mmJKJdG2DWQ1M
WUGhQqB6rc+gEKbshjMMjvI+SuawBekg1rt+ndhA9FTrnmAhDxDI/HWjFXpf0OvqH5JRv5BTSbky
j95GaytET6c2Q1GTFDl/p2bYR71dVS2To3n+o1dhMdtRy0uOhboAwl9gp1FoJuE1cd//Wu9WWth1
KrHKNlu67/fvtUxkrWl4uQon009HIzprD6sX+ZktlMOg422LkIauiHvr0HLno2oh91D3Oe4crk+g
9jXXwH5M9kdcJ9ykMsLZ/4471CqNxMpdUCnQMNwPSdOZqWF4vERchy5gT8GRO6kJ3O2SLlpQgU3m
uIE7MCIXuNI4jMuQ66AsYJgdicErKWpbB4YrRpi3Gu6TLFoZOnl3FyJaN8YfBw+5dY89pn3dl3Gl
d6EnjZ5zx0MjdrAMalPYTMJ7JyRkKA4nygB+5b6EHpXXQdN/fvt66wSOGyVKQZfWgVN1LWe3ZROj
hmps8u1tkGgVxL/ZpFy6X+m5K8wjQ0WfpyOKHBk9JcDkoCe3hdKIb5hM9hEzA7EnTtpvZQGOeo+y
LxKKpNEW56+0OC8wZLmTCgJ3Rc+HjOJK08nFyUHFkIlHe+K0ObLTeqxJuV2r+WNec2aUtLOXk5m3
VHzs7N83YUHeQIdPfQb4u1IArLQfDS8o4h4ZKwWEpxZUpCx++fmaQiBMXlce3osDvjU6AP1mDhGY
vvDpMYj31dqnExWZbqetsWq8Vlt4JBHSV+bS5N9A1hoAiOeaqfbOhiJ3mk22P8qk037YA/0wK6Gy
O7NQ4M4+NZnt3uc+cyJXPcSbKZdSUiMyMPPXsdQ/RvwkrDpUpGTbtFxlnb962zpseqGu9QO+KuKg
79MKKfbdc84RMftihUsJ9frjb0ZIGhXHH+lOwPItFLoukacma2+QOeD73S4CeqZtgShXoZKIGqeL
TULZ+jBhfZNhl5sRYysOud1habD88PYHuaGRus+5WTE6bN8fzRAxCE/0se5y2fuyGvrgZE9+St4P
V02a3srW0VuvrLpU6QI3SuOL8J2uhwKF1oqc3kPRwvJsRZdJqP2q7RJWWhZbQHyYSgXxc056LiOa
5jMRLTRohnxcAxYkLhsJiAHn2XbbPdNeRbS2X0bCtwNbDa3un3eqboHNxhd4qnDDPP2flOowjOVg
fB1HFdAx5W1vk1MUHEwSgau3bZzy+WhGBovggsQNMqLForY+8D22HpESH8h01jhs7aN047hReZWk
ni4lfI0ICal84oQRb5gsrfetzDC976S7b1hi6OJR5LzL11SaH3sxq6kdCNCRwwnLoJ4h1o4N8zA6
Hw03n4LuaCz1D/Z2RHjOMLMK8Ooh153boK3lXx5cjT5uk8HrlaQ7/v+i5s5OT3JkUK/4c0H5Vloc
GMZ5fyAhPdkeAq8H90Sl/CurmHhL/1U1HYdSb4upGYPx8d7AHINzc6J807YkQ2i0X0JfbR59Rw+A
eO1PMjPQKQle+NNyI/jPFcfHN4NncKbxr6ZQUlu2DwamoUQzodfAWIuaV2J9en4qZYzNsVx/F/7G
W98UZtCLkhNkcrxC7oqvJa1w9/A/wH94Fd7ssq7AzuP+qF2kSqF/TUjIccoOqlpCuVxUy7UfkNlf
FdPXU95++zQhFIcuMQeppD/a6KMFq5mYcKXtBruW9vD4I6NQGAdQ2KjebymwK5VNjteAL996SEYJ
+ASjZpA052Vx0Fs2Es0dli7o0p7oDYbHkOK9miTtVJwQMyDxbClATFkmK10Tk8g29aOP73QRnlWa
qcyoNfaNGWwgdeR2PybAbVY2KBFPxOUb/3CyPcftkhhq6Mp0zM5PQo83LfJUSUqcjlZKDoZ8VRCP
fslkYDXqiXILJhkiz4p0ITrbTYe4SqrU5BslR537+Q5RT2pgwESnWbCKV6Lmzo0oj0ckC7wIHWoe
qJB/J6Doi+UqtlVsNqXcZ6gfn+bpprQ6jTJL416PtavBEAdfiIhr6YK76dSib6R20Hj9pSyv0W/Y
zhQclAahKXoSHnu80MONxh/xOdGVPyz8X8aIHux2FDgJCDp0lwG2XmH9SpBwQ7jisazwGrogVQtj
iw0BmxdDjXvLPfKHse3ox1ihcXY4LdiR/9ZlbzZO8LiMkckjXi/F7Qetddkym2h+LYNUuuyYLOXT
WIFU+RUqJeZP4cwb9ioG5cp2dpNzZWbBLzjkJgc6uQlLDEvuMzuRZwoUxzlrE2jU2kgTCBCBlhSY
oqg55tJ4CPRDXN9TEmE0OYHo5UrcnamjuJXO9hKoONdtyC/OKykpvSl5QU9agSI0r29KfMfjw5BO
PN457Nr3vmDIQQlFoYccLDSNJHFAzzWLpE2/zA6ZuK3NEMLU8S7CVDvIm9DLvSRkrp/CNj58Ze+w
QwW082MBZ4Gf7MXwzhFn3iF19/hLsD7igQyfyLrrdGEY1DVcni1ipzO9H/ZTyEb0KPQ+jGy9NSh7
HoVgsY6fYZ3NU1x1zOwRLJYeivmo8Kvqiwk/hB0C9RHW5Y8jA8uu52yhC5HQovZzsXLfw7+aHzO9
LqIA6TXt8N4h5GvHcEETR1vsZC9tsUNygbaLK7JFeCLYtG30pzXfDDzTwKuEXdvQWhHYBATVacox
n3Incsu88S+KKygGG6NL/KqzYcaG87ze9AzFzNyKW6So/AmVX5XKg8fnIuNPi1UJpBQJhLGmc52Z
FClzAqe/Ubzyzo4RcrURKuJxvFHgV/yx6XHDA0nsd5RywZsyiIFrJdCcQWDSoasTJc65kYfGQg75
acDlwB6pj3btGzAfIN7PGyWP4wSeiujur9Bm7wnkgbnJUhKrr9/Jbb1x7VHBLvWEfmciZE09sBtG
Uk/TJg3AdtItfMVv7293mIPEUHsgdgkmSwTrF60qIvKmNkBCtCm3XDpI6EPMxQl1dVXYJM+WstG1
V5VYRO+nzry9BFzswXtyiR8aGBnSftKsJOf0NttwoapFY9Ux6JwEmERrMpsHPELFaUHNWDwm6QOe
fwtlIFP5wcT57zwCZ8jpqFsEvY+ym201VAyvMxYsEYGY3rscyKDHMJu/eRvrRR6stGbSpFLoxFtZ
HQVut3kMQBqdiCXqpO9numvGkOhvQ9O6jOPapcH9RbqeWUZPKzldEKQTilg1+N/q8pbGyqkYd2Ad
Y+no+TrkOIOu3KbCZ9tySHSbztR+GchCWLz76jRDxmxnhSC9+rW3m9mAA5twhnfD+BAF2hCXbxnP
9/4r2vyVbrVTf4nF2SZGrsQkicZu2Mcbq8Ajb6lk++GqJfnMy6+lMtAegYD7jJ8zrckR/M22jl27
xSlSx4FDU3Jmbp5BY+Qi19d6TSV0BWQVCLk4odSwKjzdv2IWcVmUuLYvXJXw/GXJU4EALxf0j5gg
gUpWpdUl8ZqVz8jXbZBe4QG2Xu2gj9SabeDYn4DGYfhUJ3uCjbeUO0fDxezj5ezDA9ewqDmaqogo
Ull8dgNc3+/LcnFaEyeyODIiRrGTZXe48wHB9Crd2ysfS7YBTeK+B3ka3CKRc5flb7ReVCXQp8Hw
+Yk8/TySR0IFnc/AmhQFCdPz9/RvfMmVEulSg77t4w9IvXAs+bLcURz17xsqHm0TNzRnf//gUb12
Zj+gN0/Gvy1mnXhbokBxtqh/vrc9iVKyi+unfLg370ghq7ZXSSy2mVadl161BIXfQ8g/OX13LiO/
Kqip7Zz9oPfO96ubNa0QCoOjEtsUTnTYi/4o/dhleXMHdT2X6nJ3ehdFZel3dsYwyuYefjqas99h
U4YetxGxxljSe5ZsT0O4ULr90AoVIz5JrZ6EYKPXjboR3+sVJf5PLHiIbggvTe0pg3IeUVCb3+Bp
V+s2fs6ukgpn42ZzqCyE1wUxd+OEspU6N7BTJ6Odu0MVIKZtETZG5UvMzBs5BOhp+YbD4KEmJagW
zPOWzQtXrhoHZVkMcRnaY9uBvb/cMKSTwIFgwuXvK9KtWbvdQC+0dtIGUetUmTgd+N9JO29IK/1q
TW9kqN73+qJtOLaVMeniZmoyqggv469i/JycCi+dg/iYChUmQPaAIFmaWdoqCKToJtxmdoFhuc3V
NIFccl05/q2PtxQoLtw5FBLGnkrT9HLdcH62qnCXTodKC96Og0+6wtIGyvddmdaGorbSkqYKfEIx
3VRQETpDN5YJ0YRpL0QUDh3xSHTw3rAqIApZjof+O5TwejPFAQhV05FdtM9OG8ua/fK+VTF4rtnS
VIwknFiZA6z0ERyikcQSYdLhgiUmbS+F+W5ArMRjgqStaBeX5WAeNCDWPNcphq2SXeFdsxOXTV8v
WuVG1EK4mCMP07Eq/0QkEhMAMl9pmywNAwbvNC9g1G1d6aSea62pRTHq6sW2AOuayslmY35X8TCR
fpbtTTYbbagN+o4LkfR+/ftJc3GrwZJhfXox1uM7Ad6SXzo8o3hFoMuFaNXu0Fgz7AiYcScQ0jgu
k4T0kOYMSdYyKJovXmI+Y7XinUIZydXbvuWPD66jEWf1tKDQShpBmbo4rieAOENKfYFxBIsowOT2
sFHHmo742SQcbgkgyg/NM+fR6fyivXv7kTAfffMDZQPiL5ivVSURnmGQY61xZPDJivRUbS4cGWnh
fpBGuRzbcDI6lHIm7t7kdl6uf2L+ljMqTT28DZnBJQGnu6eaEV3LgGI6U+hV3eZ9wc+uBFte228h
Xy2TTslWXtas/H9q2Y7Zw/+ueho6HpxH43CH3icT4O1kqR8fzdyb6GivwKg5WMGtNz/MxzWskXP9
jMqroaJ3Nos/mrsio9tf+CiQr23dZtNvil1Mfw5rShmH5jVPazXlNUoH/qWoWuNolIWnWDFuzkDc
g4vkrY2DBKmKcq1jWtQGC9MPjsIbuSCEKnvkvZN6ODbmuQe8a5z04SvkY0uDNgCMg0Rb50gRNHJN
k/lwdOcdKBh2piqvoZnA85jyjh5li7rDXD6MbJpKvIYjFhFZvFYo8qxVoUmGdSWkxnrgvamELjRm
O9f97bbSyXRhTT0JxnnMRF0pPvz4A5HFb7xryaqYVhtrQbeJuHwCWDb9sSI02eY21MqO/rsCIBTb
r2nu0gf1/at6ezFVnkOKFNiyNHDMrJJMg0G5ffPdoOldfPXP0SE7oV8/odNuGlKx4i+K81IJQIsb
j+lJoGjPrRhPGKUT78lNj0WTY6EVrDEhOvDWzVyqiRDnkK5daaVyfsMdzSiuXmKnUObjoWj3alfn
EpM4St49QLSaxqS4Ge22St3NehX8aH2XIJCADqRyRHts7XkIanT76l6Q+pLuqT740bgGymbfVXOV
It8O5FputX2dF5XZBgaWFkDuOpUzAlAalGmXpHpf8/UFFGNPf1jhYxDwi296hEmae4X7Ajjzs5OE
A8bB+0Vwh+RWVcpZPIzYCU+PlMOTltNZsU8emhrAUL+//yppTyI7g6rurnn9EDX3+0u8gZDXGMsV
LKqIlP95MrAZInhWEB+WSmcTtVU0z7AITkH9VmDhFHpqobDTUkssvFPCUKgKsWEI7tCtn/Xe1f/x
1goBk9kfjViskKlfIRdulds2XUpzJ9o/6xN/ZQGlPI4/Y80D0gQZ+bfzbwyKKI0cFOpuPRZk9/TT
cXdYFinJ2VQEdw5NPmnRx/+5rlnUzLOKDr8xi7I6oAVYNoAzsy8TbFmcNituyc7BI6+bwfQvOYNB
ldGi/pmocwVxccRy4U6mB3Bid/ocgqXmkIgUAnvEgyZCD7I/JhOp8/rsIIdzgu6ht+1MEIPYOdaK
7V5E/JcqiJ546ur+4J5HfYyyciaHIXwOsttEgQOyMeJx53FIfsuTBIxBtu1ugovMhrAUI3BBB8fh
RLKS7KoPBNZ9QTI9UyvuOzABoENY7DAuuc/nWkA4Awix+JFh8Cr0n5ziZTbpOc8J9EhYtKLbJ+85
oIb6V6Tu7EL49P3iuxNBUMGGSL6v6wlRpU8tYb9DCbwpjdnzl/rU12a5FBnBNu4XLKhIAjOn2aBf
uROTo9/dKBHzRQ7ZygD4ZsFAnB/+4Ddp/YW9U440LqaPuW0zML0Q5lN5PdNC83helASX11d2l31K
o+zHdDJOANCN+qlk1mnRvV62KJ2GX5XmFQoyUyPM77GOo3J8RUeOjAznTAPZFzwwFcqgmb/8C8jL
wazzOs2kiqGNptpdLeIuwuhU0v5R0PX9ppBhO2N9frwISgyUc0e2dx+1atIb+7wRwW20G5RlfD2/
JK5LnQOXiAPhnl9lKA3HQuBBR2DCceVgd7caP5Ggz2Nq8TaCEjdp+OqcGPFyVK8BoTjj5s6ST6vx
D370WsVQxfnqQIu9U56oxdfdUHomekY7vpEjPXgJjxQ+TbygwKVXcnaUYesgT6Ijms8c1dpk588E
Qi9AOaRuL2LGUngmTqcQbtRJdlHm4DE0vu3NJoYKLk6cj+k8498ap6W63hJE68TN8TURxJ1bDspN
fvKunNUr6f2x3Kefk9x+tov/X1RJg3PDg1urIYq6r+WAMS6mjIcbGMcfYnLQZYi0MPAGEF3kRi0q
kHOciZFDxT4H8AT+zxZAMgWqf1+G1bstdeuZB273lD/NxzZFIXI0EYQewWyMr54VXdO81LnuSHvF
QuGstntkIoxRXE2GlL5lV1cKkXunRlkMRwItdfKInOdlaI8CyNnq7e/Td8IQYoeQP+mu3cUw3jK8
Hs6mJ1H0LSGF/ykKuYUxvp39//chKWzQrodd1XkuZxz15o8SrPtF1IvQG7X4YHilOyRNhEtV4wBv
Imxc/0WrJUkAG3HZ7j9pVLOP1fUwvfEeATQF5wp0f+qHjpdhrmoqTpK/Gj80qt0w085NgTDG/3qF
X/wPY2N48meog74C5hnRTuuutBvTFqRM4EdRZj+yLjg5hu54J0KlTd9hnR4yhU3bfdFHZz1U4JgN
KQhOmWgSjwoHPqE+bs3168JnSBS7BWiB8uJqMPOmEHBRgVuL6brycePUeDiGrVrVIzwzfwUxErC0
2r95Wz4SjhFX8JDehtqjQaTcNlCRjku7vwXqIUikcWayivTW4zEuDLWMARpwSPDG/FsYVgXUHzGc
8krYs+11HRS0dKJxc4XXwIuFdG3HNjTtBmZYJGCbvBLSwrVTmf616fBtopI2UNW7YTbkEqR8vmhl
GaVF0sLH3j+ZyoPJ4AgtowIgVEbm9XpkkhmPjhXkVU10uOY+4FbeYfGify/362KvxQPVjbvPt6KY
HsaJRYC9bCMYCoqMr6B5I+ryKNwlGUiJ95HUomhv8jaM8VI/bVcwq1F3p6YKKrJ62300ID2Bbulr
BIuOcR5HhM89+5SXAIRtDDLPGuuvKzbnuaP60lYGAK5GzhlRnbxZFLvtjDQZtHoljTdi56sZwTEn
kThHma99WAKyzV79ElKV/zlyShN2AsCTjXd56RS73VPlxBo/3kZ35NXkUuKxYQqE+851LhL/2dHO
MCvCLXo87233mOeGpQP/AoJTb6qcj6jIJ+ganhiYoOU6XY/IXmwQbr0novFK0PYLB+LYS+1qwWYb
Dh9ByVqrh47Ll3GYNlKHgfagXeuyA1Cm1/rDyja4rIWpT1IS5fE3dIbkEpZOSzoyZQ4a1IwHDrmH
2YH5jqgLYBqzDEg/l6wXFEqIXd2LTv++IgTkGLrHsLYHogBTQDF/0tWY4Rw2feQ6GNNO0jh37tbr
xkEshXPuuY6kO0c/vO/lO8JPShj+EKtBSZ8c+xJNprkKadAdbfUEC9pyWz/oWejD+Qnfsi+Q/FQU
osLRFsuMSnccT0wh96h4OB+MfYbdLU/jyHS1ZAKSjagxPdHLQcL1vwM1QGFa1RKur80fT4X93nae
4lXU5K0B6381QBM9z9+dO+vxi/f3yudJlrHj3x+9fZ58gro+fmRSFrCMa/wxXJVgALAiPf8ldA8O
Ri/Lrmwjoon22oCiTtJDjpHRs5NWWgdmCppdqItsVTCTJVj4BH8rTeTjSx5bt8OmwnkUO9xzjw3V
hI3QqaQLgHwvoKpd/Pgw8As24+dpy7n3XafP8V4S92VdrUNKT2CFq4E89E54s/6pQ5hGSGAJ/CyM
bYXsYUn6XU6u+vtFmxMxW0Lz6IkHe6ujMua7oJt2SThYbUD3CjqwdzzTP6eo6+h57UIF6Oly8mMr
UNq+wzhmkPQ9ZfPTuHPsD737odfHINaz6G+Yno+7o+9hyihlXiV5SwR1qiOO7O2yaBIP5kNLfqfB
OOxmIkAdVRh/0e3pG+jcCYM1h3llk4orBK3bIA2WT7xjUszTDCIUD1o0NTW2WhukC0VPTCZUeCTa
RcLyrp7F+4+TZ/HsQiWKXpo5D15Jdf1HQrUHm+6QRm6uUFvhBWGLc9pFC8z1LT8GvtOfM5elUg0d
eW6InR+qYBp+/RFCs2U/McXGlIxSDAwNzcQj+RsSQoYhzQ78QZQm759N09I7ZR/jObsg2sZZ6sBb
1tEuApRFxFUMADhRMtEhn5yuUFwQVr+k+n0ojyqhn+DAH0Ya5EuAE6UgRVN/5TrGX+MXabrtX7M8
0ea/pzEcMyd/VZW1+RfNj1+cHxj2gHXv3H7rIviDrTdK3zDcS0ae/dASCFFMW50FIZjQNe64ZVFw
Kt1NQMVAwf7/rRgVFyS4qNrMuCqmFK7KIsDhXtzTGzvuTCbOkSph96Mcwtfq68YfCXT5MqqIIWb6
h3IctLJiqIvLzcNAtKWMUlsgSR/msPjhI+NYrKB+Yo+qpNOOlFK1L9pimQArCzuL5fucisqa8X+B
Fyb2RQygz3CCiI28BFkPuL4VoY5rBzFF3YE9jDsktLkb0pdUAjm5MoFnZi/XBbyQM/GJ8TD4HDN2
BNSBxhtvKNMqJMqAGdiyd8hopbkL+vVuSG64tzYXe+gqfVxMYUR+i1iEelce+u2pKHEFH6qqkhDC
tbsgyeH3b3Typ+csB5/+U+8AkUJ9zIazYmuzXWA0nofphJmRmTdYIcWMmGaYXp3FU6OzP3MmvZwd
cU8p8rUwLh6U/jcUn+p1zJNSqRDjMsPtLghel8V4uE3/PsAcS17EqiciE25zwSx9gO81iS+D5oeG
MpEA2Y1raoRAyCzYxxNZgp9Ng/Jh3ei0pe4TNvUWetudhaPIDp8Vh5vzrnHmX35XtTJMhoSRERNP
qrwl9v+FSrFoTJ80oE9oem91IiBBsKAR8SNBQkB0LZB0bkYFi+SuR34Kw28vmvzHIOuJDzzpW3Ay
sG/Nmj3uJiVpUSHxnpzMeziGy+C4TWzXQt1FcEdEoE2rPu0S2iateMHP2/auqTyfno/Xx2Fr9HGL
RT2ooLIkK+T9sAV58Rw4arKI3rXTxSOtPzN2dqTjnfIMnwASX7bIfzbmf5vCRvY0jrXxg2WcQN1p
HBebDgr/Sfj17Vy/3jMVMLYrDrwbkBDh/xt9PDeG2O0czVTFIjWzngb3BpCZUz5NdJCcB42Q9lGY
41IMxLxupzTghCUGOIm1eN4OTGDIHhvCcF3rZtMiKs8vLW9B6N5mUd9z8iSkcTQ3rXsrkQFbDdzm
q0DHQexozl6TiyhkWOQkqMetYtyGVowN8kBNpB9T5YUmk1Gee8i/0KdIfapVIxijsUDb3sVf2M3q
Z3ZdTCWe/I13VCNW6HfSfRsTKoHkHRGsbgX0SrloieUnhOKjvCrVx9rW74xx8BOoj4S+UDJOSLFr
pCvZcemSJpGcjOOT3OUvmeDQuw1rajFElgxkgqyR/UGdqenLfEzZBjj+6jolnJfY2JJZiFevp8y/
L29KMpumushqp0DcfrcfSluZIViNAn9JwstWEbWccwdJ5cumoJOEMn/Xm72BgZrBgtwl3CwCENBY
oRSKVeR7p8SZRglTnzNAbJq2KpoZO9Cg0O3z1mCzZCC3arE4ZkqQk4ZeCF4bBNdKg7LTau4+JJQI
AsxrODelT1dmzCGVQxMs9s+uOQtAx4dQtcptGuOxsu7EROYcWnqbv3wzMmGYXsK1gpf7bxR+880i
j6bI9CnDPUCEWS/LWsFUYfyymQrTm8Bjiad9lQ8PtkEct4c6clGWKV+QCbDH+wh6lQ0fCPJTkMHs
HIWknWtM2QeOcj2qgzWDNMHJkBsjxoxXmsfF+Wk2bu1ktXe9NtGt7cA3vpQvy4CIixoQTgZvP5sy
1xuwbPDbdk1sBcEYL23Ducc8+I6mN720DHfgC3jBWIOOpg3xQ/kUKdP/5FK1SAxZC+XbKTX0iIYX
iWIAOIU3ztRJXnKc6CBfi/Q8kyG+TVKM+jkrD8OzcF7YK6zunX7kYilbEpA1eV37BNP6NAQTTB9p
QEedU3+/XhrmVoOwaTkSfgogsXYl1YMxk8M1ghCr7NdODm0DczgfClpWg4W0iAnvMWpd03e5dHu8
YA/kKtYo2QHR2ytW0A9wGN4bSHHgk0T0wbVzbf6egl1lH5O7gs4GZnqveR21x/sbf8bguIx8m6iF
yVardTkYzv4YdiHoJiqja5qlPWHtJjHP0w/M9KySOm+XmYwmktQfFwalHjo0Pozwv4xo/5rAvPad
b7ReyJVPSW0roE65xzxj6Zn5YubcQy8SAYKcapT1nGU3xgbNYcLHhbz2d8G8TDkd8C0nkQsGmvS7
GYsOX3W22H0UYLN1cmssfXoWk81TUfJUOV281u3Vm2y7Mtqm5hl/d637X0naJc+BAHgj1bzQJN+B
lhYpx68fQrBztjSnY8qIva7S/0jU94FwRlOcwOGDz6mivzz4LsnAuGn/0PfVLTy65qoAbIwLeHKg
mSeFkI1C+KF+gsZPYGvOEmxBhjrYvej3ExAn9TBhp1MVPWNh5pkh5CuuqtN7iwvL7dUEmxudUdUs
nbfdSdtu2yVH8EvNFdc6T7oUT9SD5Tvmx1tz+7HdRtYCEIfN9/CGcBUyBdmepEx7bqprLayeveb1
mnmP4wb7C5HWFwX5LSUfvJvj+ka5yKxF89PA6D0C4St2FdZTlYuFH9UF0KvatS/HvMhSWrFNwx4G
lU3nN0BsR/La/OjstWeSQteBQng6GKIdOzmPFAn5HwQpQTAjmd8waErE+MwwROrFbhR5zNeUhZZ6
pPk0CDQzqMOKaUdq93vd7b+J0OZq02jey6JOlgGBuW4X4aHbJPDcGLMEK75JygIzIRXUj0CAgNk9
dq1GchdCBtlUmGHJxGI0rlEhr5r2UnNcQOa19pZxx1OYwjM6MPxWP+MydesVvPD/CXGBR/pjEJNI
Ps5VGJJ9JxTjpbth3cBkB89TZc6kwZ9SpU81q5VCxkw3yMYhVqy6dRBs5u68Ln871D+fzjMyzpUf
fYYDRXVoqEwHCBeebed1CpHWsayzKPyufojsrcHvFJo3I60uHuQefjWzXDn/5J0ldYIVt95ql/vw
0pV2dvHMa+EtVODmKtf9PgmBYQ1TmrmLhM8us332UXPdxhi10rKP/WYUzIAnXLr5WSqex9mgki2B
58ESQz6xQBsvHWtfYNhvh27AxIV0SXfg1/x0aUzHDNcxQsbYwRCwvYEESKoZWP/MwwXMgTAO5SZ6
8eIlggY4mJrgUYk0NBcEtuD2VQdKT3230xL1YgR0KIFzS0N2a4D5OaMhCr27v1OD5WLVjjRewBWq
WoLMr2SGsyxH5Dzl6KBA09F3ycMBcf4U0ECOMO3yP8Xhbsup0eZ4o1jTHz6zfFvZz7wPsz7AppUj
91+Eg/4lS/M7ZKirCF+1PjPyxo+jTLb+irKbloqfwSUJZhlAmThtJ/4ZVGotWm8VQbxd4CnCOVKQ
VuGm2n5UbIIeekj4dBhYGk8YbZpK7NnbBHcpz9x8NNlKzxT/t76ikPwPrBvw4n0w43KUGyCFYxJu
d+7zIJsqwTGAlvI0Z1605ZOnvsbiZVH6Gbw7ohbvBtEwFeDmJtgEwSb6JJ4mlB2M/WeGsj7w0GfM
FDjkXipDE/gRRVzoqAU5Hclo9Al4IVY9enE45NW+9RffoAyXahPsgby5g9Q0k2VtBi25tI4ZRxFG
dBjhNOkZr3hmer9wvIjoOsa5yaUCDlvi0yn6JTubyxSDgu1mu/WE2GHW5A2A/OwT/Hi9Ff5OXsKP
o4WvDmzE+/TXQ/Mt3OfiYSex8A/bag9U9JQk9/53B5l8XzYx2ntR0Qm+qLe6g2rR0CgN/ovAjXPW
sRe7yXBhHBlXTFEpQ5shWwQANHl8LPdqYeChWaDMi+DHkKaiAZKBpHMu8LgQqVqfkFp/m2AR/nY7
Ei5SS02nk7E0vWJinWqv+r9FLcbsjHL/K4s7hfKLynHU/POmalA5Hm2+EOnMuQnQ4ow2nKXafEAE
e4ZRQOKR22iqOhhodO3fqKp7bdDM8dH2dSCqAi184JqUF10vZbLoH1sXmKZFU+HvA5nQma7V6w0P
EvglD/fuUYWrO5yY4nlTM4BL+zrnBj6c0ZwTKxpbNgHH4WotV6e6oyCkwgRIv4QyCaA7H5xiaELD
Ds8/4bw4TZLo38qR1OIBP7IieAxdqKaTtd/Z14dzJmRmzt17Cs3qLJI1eDTTjFTY0A6bR/fzNZ9l
gYwpYPbv+4X1ulbdm72D3CVJYXctolu/7LAZ5AjekOPlQajCRmdoUwLH0Br2OGR1w6fCu5OU61hM
+xtIm22dCvTqP+Qhf59Dag4lMVl02r6NPW5S/hhPGTkppYUpwlTjzYGOuajZKyO6uJJ1Oj1cq6VX
gYRSwVGluaEKFIS90/TKamZDVBQZOuF5HXYn10qKEhinvvu3UIg3epjHb0LWeAD6wubW8c4Xoh6X
bniwSDpGw7Zhw1Gv165zZpmdA+CG9gDB9WFnMRnvPy9b1uqkB7Ps4wTpRZ5q59LyeqNKkVn9Tdto
yZ+rxk8SPNDnLZzvCPrpTWbMxmzwUgU+Q7sI50oSAbQX0eV8voFqlgvzh2pRwYtmsUENTTCT9o9y
7kyLDAEM7KXN+lrUV7t2zrfM+JVWo4NN+x+XGMI+5BSbGLQK+CgDekUFzXJlddqKOcxvEYHYVafi
lhWQAmqS9v88TXuuigHT4vZc/shqY5B9g3WqgV5v0ReBzaWj7X37yqc0Pdu+4XXihtRQTsY08xii
RCSGdLqpg2+p3fGqRQC2IcgN4T0W5Nrcdgs9WE9bKcds1q0VUESNM6h1j2d+YHikon/tQKvFXnam
m8JCUjcnGsj+qCaXCGeCqmpiMe+LQrc/gy8JnFxidOXzs0Tm0KLdbwr9aVRRQvHUZ7oC/ZP1Cjc4
tGW7pUhFrATrozvskQrnqc0Vi++Dsu2Z4eX7mZTtFVdYn4mxcWYbN9OA8XS6h7tvdYUzt1XtM6z8
UMS6rCdjEQgvhUXHxIWFtJeEZuPEik44QMI+9snsn+N3xZ3ptrtLPwPJ4aVGRdyhcg7EFz1hQOu+
dSlYlQRnQJSU5lQ8OzbFI4XcoN8p/9V9pjoLYmbsALieBowyHYqntl84ChTArG6PM96ZrPVREZAW
mkyqn0V1vs5ShH4RrCOk4IEwC5Y0PsKtPh1jcjTp0Le2UhO7iMVX2irJMn2Giba9h0FK4NXqJpaj
xaoe/hfQuGEoOUfUfNtUQM5wLimKACX89PunCDd6Qav2+Q1oUUGClzRdQoReEfSrsryrUbNGApU8
L6weVvoUfiLvyS/Bu3gGZ9caWfAaTlh/RNdwEPwRJMgO2WhUSSZo3aF/v1MU+5CcIcyMDeo8HBzn
m6OMS9wMgu41EurXcueYWtsV8yi5ganhmbvEFJJgmw0WYHsZH17iM20WulA+AUDV4SJtGuO5F3a3
7x7fwGeyEOEdVY8b688n4PqtXxo2KHLIJGfqrHUwLisxYfDbc9YMGWiccKVxUjLvDlBQ+NzhYuiY
HNPVansftPtpxl9XybGJ1mOlky6C2VWjlozVH1QkU1f3NHJGJkphqm75V6bgZxtQzST0J1LSdDR4
Qu5GYKN+Bq+McQp2loxAH2AlOLXdneZGULvRm1q8e4XCBdQWWPeBYYCjKLc/T2REnN3DgKrUI0rq
oWS4QCYrvhWLYpqUQoPyEKKkLj4zLPBj6qx52x0qdTLd1gyUOKXM4MgaxAKhcSzW+cNU1wdD1t1X
fbu+tu2jweuOlOUofngsUbiPNlEhC4CSjE0+Qj2L+k7Zw3goeHOiSyrEY7ninMNvHboxFO1qlGXe
JqXBybqYeFIKHcEvYbjPQs5GfQR4dq4DluhEl6GFN+ZZw3EmmR9bBIs0mmEqMLqb4onGJ9cwEqu5
zpFKbqvPZ6TslLn77HRgqfQ70nimgmqjWyVbs4tAN7ptBc3KRwTVA3s6vf0IBKbTqsXCMA6aHajB
UNm3lm5vCqxBmkTX2vNPbtzW6lDisC+oUK2n/TynkMdZ/zANZjBHWmiTtFjPqcDL0+c1rZJOhOUe
O0V7pFVAxA1OJGGvT0OV+6SUSAJVQN8c/27ApPmJ5BS6Vj8QzJMylaHejcPr7+LXyztheUF0xem4
cBG81BnH4H3ORhbGnYsuwFtQlJlqNhcpGTPgUUUQHPASr/J4Xm1OgKU6qx/WQsUqThtKTIkFRxCM
XIIsXYuoZTlZYcOyzfBuaWiSH39VEiRUc/yiBToJbACO4Wr4uYNjCoBOB7D89eG9VUZ7H+cZASw3
zxUNXPl5BbLlz3vBBjxs9bHaeHzEGn46p3DqzrsyJGChbIMstVBE32csLPnHygEHMr0OC/ySexSd
Y6ToP5ljz03KEztFQgPM8ALlBFpy3bJJfp15f724nRGFQ3rD59wrJTtlEL4X+ZmCLD1fcJLSJz1k
cSBOmiKow/lX4kWlK2Qqy9HYoYhtMT4eM2DxQdRpR4Z2ynw3CMJG6lgyoBGuDmcryY2vDomoYy+A
djo3Z6jMhs4iE/EWBlyZPThVi/zIT3WHbvw6Ow06//DfEKIwz7O2/A+Qes1PNwPOZD2A09Bmhv/A
bREem43LppZYmTSpm0yK5TnQdXCr3nW4FZnPMSU/U67mNLkClv6HFnakR6ftMFCNrAAIXwmJVR0j
4/MqIA47S8A9C9YBa/k+VYzd42H70+SlKrYFPOAsTjoZJwaXh5P81BNi6JTrF+U3m++3M8jgyeMv
z95V+TdCwvCjGAfDLXrSJTGAfJT9kXd6ITlfbZ7bFE0Z/iZags6cQZIXVCDzaOTuGbEVKePyeJJi
fLLaKvSjpKMB+XsxZpfbLhTtHRB207RTCDroibRLcvtptqxoYaRdRQMFgKwlSO+zGYiPeUWiGOV0
WOk8K7cUcKfzKvp2FqgHbux8LLdbGC7/0A+YwunjKcAdryJLHaqZU5tuMs8czs9obSm5fbeBDIUl
OQnDlZRvB3S14VmXmDpNJagD+CjBtS8oy6waFUoIqxgTEFJEOYDZPAJPdT5vFk/powCw5evPkZg7
gq8V0Rbg/vz4uHTpd5ZzZKYpz+/pHLZGNTxtfZPNT5TBulW49pUbF7tSf9pFUTADZz4P7oE1qyEP
M2OpQwzgSmT6jZKSOmzzK8UJ2gF7SFnAiOgL8jDZhzFJck1v1GQB+Q4+rAkQgRnCqtxXNLwSrgsp
2Kd9L24TYqJ+kdCeLmQFWjp+VuEBQIZ69lpNxRaXeole/75qg1etn2tzlU5CsT0mcRv88revHQga
8XjanwvlML5DZiNNNTlwZCGv63NUT+cvv7IdGBMKSCDgmetVxidUpEWY+s2cgaQZ0ho5efqTft6A
/80KE6Xj0LyOCo7RF4g8vH/49XQ7WccMiMDlZjnQMAsJ6STbKhBJhwxwEO4YU72PKGYPviyk6UQu
/drYdcOkxxQLTDz/JTZ+Q6s1+7apOZ+Q2BDG/lVhENyZDLn2vcSMPzzO2Pub805koQvZROTb6Tav
EqC+L2KNR43bW/YFIftpyLJCW2A03Cd2wuEuqhUgGtPNVibMYVxIiagTMl+MPC+6wfY8M9MD/y4Z
AlQ/oLCQP4U89Az5KR4Nov2fwePbZ5kR/n7k/7UQq0u3fmHeI0e69C506MMXttNCjZ8F6oQclAju
vOWDgQAaeHfpdZhTLMK7yqLvosgumS+Zg+fhydYaOvmTUG4R3awNBhlBmkIy68iIKOMmk0ku8s/N
SfnIpWDGX4lNxinusY8NpXS1yHocbouu7TCwtUtRAu1MCDh89DN+iXQLf6wLQTudDzIYqLG4N4Dw
YHGBKxsNXjGj5ht8jmgss65lFoDm2Od0wT0MT+SYzHQ4oKlccwn9ARmvy1MF3mZgUuYmjmIB6E+s
bE//iUOQBzpj2Tb8EguLMflXDIpSv0osiwvvcRi2F0AfEvdjJmh+JNYbAAPL2OZQCvmxOyg2StZy
L0rGKcZhr7ynTBfxkba1wt8KMJ+pooJGYeNGkUrT2oH72qMLuoSlBNYvg8R3/pTruUrXySjc/VhQ
+ZAJYeNuOGguL+F6Gquq+h82yIHQhlJe27hOXbrBfkyXCVxPZoYSztrm635Nz5N1t3+HmPS+crXH
C23Kl5tNY8fLiI2HikBdzAIyyEukr21XFj7rpO/g+RQqOlDURL1d2VuH6eyZjGRUUtLAmW3Sbk8d
eIhh62HQ5C3gPNcPz5c9z2NaLpqn4GaORHM7NTmXJogmHWR+j4l9UL8o13cY/i4uQVwFc8fZNgXl
YFNu6izjtSUQoElIZsFz0r/A6TU6XZAArtrVssutJF+K1PzYanEqT7hEcK1q1+V+KnAeTmov7PNJ
eB3855J5HZKyBqEYgAKQQG8zM8RZOYZyFfISNn9Hr8G3Ck44JYrBXIDN7vv9JDQTIeiTZ1jwmH6e
bPnwMPp/i9eZf28/D3eHhR013l8DKwz0BtoYq4s5Lla+wTxMbsPsBKf/6cDOKtVgabpiuWzCI1YI
cx5Ge/eBHCkTE97QIiAL2sofDMl3S7h8PDPWaQbDH682wMEXyr+ueMnFBX238JN5KcaMsiKTlvnA
u0tdjpbCxmH5zuF3qyr/EWUCUdwR3K8+r6Eayh109gklIwwupO9S3t+IP8N3LQb/G2LIeFtjG59U
4C92dIzkbC1+w9w/iMtA1ueUBePPQMnylgf8DO2rIhE195Qf+b60U6MJpkuzUajViegyqNvvG94i
mx8NbPFEHA4ZeYt6ViveZBG7LJ1DyL+mCuf3JAw13Dwdz+cmmwAuRW2IBS2H77WWyHHJP1Ztvu+G
VLMTkirpP2F0EE04/l2SHK0ByI7W+POmxTQ/eh1WfMO8HGXjhV+PXTQl36EuFPAeVHz1KnDFUI+a
dkZiJJf3J5Mk8oPkivragUbW0stYKqqx9O0ioiytT2LP8+dWyRUBWC7Hlu021Dsya8fhYL8hLFup
mF81UrAnauC4RZMOnsJtd51LOI0kij66vw64QlpE9WqCeMsBu1CJriHR+ZPV48mLNj0AFk1Nzda5
ZeXd3W+gDaYxD4ZOEdVp4i2zu8Jj3cW5NScoE//J/AiWcfzd3MNQEtrW/Tmktpgv84PLymk9BOCS
cPV+2cyat5b6roF5oposR6qnOMg4NaNEJ57BKKXIYeb9Ma9xXYLeLZ7DlensG+K46h6xjyp7SWmm
iap31cHI6JXXXIo6mz72Be1bDjvM6saixkOL4xBop2sLGOOMe6hDSo+YfMcvdjzEKSBVjNDnkxkS
VViehzgvaF2k6IKGK/rcD0DHy67gDe0n0T4vdMTwHoz3uZ5P3hGkwxslVeN0t6E18+6K7/OC1ZOJ
s71XgROVyMtvF4++EYVGT7KJluCdkkWC1YEWDnysuw39EkK+SVNEYhsR59Uk7LZ3nHk39MqwKVVQ
3iyr3qNdMJs/XrxOwlBXaGInvH01olvcF+Cb5VJczZtHqHmiWu60wQMpTHrpsltir9tiYV3mhUCi
P2gYxoEC8e2WzN5XK0GYhEwRqZr6TuyzPwjf1eqwKKrkB7bLNwPV6KBwGZI7TeF+92M5ZfBiwI9o
JejWsElXFYdOkso35eXhfMUx6+lF/c4ltzTblPeHvZoZJ8jwHNlXXkALlaiZecS42pHW0Msq3ETv
e1f8tw1vgduz0MNtJsuuizhnAeKSdN7kgeYdYaHE18KOMeBX2fK52rg2V8pSfAvPR8NNnItXTDBY
q8d1sWwNY0w1pjBcWpFu9TaDuLtOsQ50+yJSVxy79b/aP6YfDnXELivGHu4ESkHrAzq9jPqaKemU
0H11/RniQ08iBhp/QqaU2DiOYUidt2wmlzcXXpe7WMKeNJzP/5O09JvwajzMkBP8JOcBnXxR7nl6
9+BFkwQyGO7/u92s3yT4GioaVNcc7gH7INr+JazAWX5YVSba1K3P6+RdpxXZ9tAn+EcPoqsN2UGW
rnBA5B32Iq3DivLPW3NAYcMK6vxcS6sT36M2rJaZ81MQdJYY6C9YLbqeXovIwveX4QbacDPSXHap
epBGDvM15yM6ZykK4wLNwIk6EnEG8UoOYJ6Yj6H51HkgxteLaL82jv12ZlmOX0CWEFyLG1UgNpp9
H1t3K4X7baTPeYlHKE6Emot1ybvYpXb1RFvW8HDtf6BA1GaiXrC1uFy1tg4E3q5uPZepfUtfUHEk
BGMbtsb7SpZBqNr8lUpCdwH5wNgv9ViWaBHbXU5ze19wJXQq6Vr5EunD3aaDaMBbFN9CJfLVR/uw
fMejeuTIx7xhD5PFbrTXYmNWn8J6I428jOML3Nfvr3G3MP7CaEYcv8XC0tq+Rpdn6nNJ2GjKRnCH
Jj6pneQ4o/wShfzfuv6+8TEaZImlylyRhcZoobI9LTmP0XVU3uzEu5aXEBlXLPV0EnhNpwxH48HR
sqDlDi4EvH9znwlcd9pw4A62LyJC5mjfkvTvxbp0rhEnT13O/ed51C6ouyImB4ajusWSRYfuE8HC
dXDkMGvekldjXa3kcsmCUW0loFL3u3X2wCdDGm62DVZr0DTJL2qnJi9cVT5smS4UhEbUwV7EB6Hr
QRD1cFE5p+3ai0i/2rnchS80XOX74Tm9qn75Rjzo7Dqi60Q4FbR4TFYK/TQOZ7cb9iog7xORpudD
gBm/vHGTGk3O5xdWkWK+Q6qpLXtig1IKOdA5aKrmUWQVla1Hna3N+g7qgYSFJSMQvvPOt8eg22hr
QC0BKudTc2PWanFTBZ9AMdKGzu+VwzCrvOWIj4MqiQ4eDef18FwdFg53a16GdyuGb7YlDvWwIK5w
m9B7HJzvzELiOFW8AUmTUIWmWACZ4VSqXJDjacdmcWD80awpx4m/2Sm+CsQOa5piS1sFpwhJeD8R
dOJXyWQ+DECaQefIKUanJOBsAhGzwsOPebx7VobOFf35HMvyqNfsF1t5Aelh8iM4uW4cswjv9JQT
DnOP4K1woBM9TTdnymwXHth2rF5UNxXkYVgM4gWE0lXDbypGreBbC+aPfNMQZOEPbe7jsMnvluEc
fyS0g2cqFc/G1zih7pLuDMoN2C7zl2TCwe4x5C2i6TJgDB4dNn1UXDfOMr2K506vjLr4LiaE5wVG
YHbiBlqJaC186i5XzlDcLllUW1IWnCBAzcaaEUugyo4iLwIBCDZ1WZHRE9uLCDotYcWsXm+N09Ih
62sK57cfR85C1V1iVxzbSPUU7LiVr1yZqvm4jpCn0uJ1RC1pCP5lNO6HAV0U0Sft72gSN8pcUFhf
cL4FXqDrSCG0NVfCddfKiIuf3GHpmFBlG9J5qowzYmjaxS1QpfLJieCsFjI4nKULeIoHGtBsjnUL
uy+gqSInULrSYkc8NW3//DONryrv5R92Axs69CGHFcL1qChgKSAakA6vxfA1xfvZr87ucG+nyg0i
SEnCyAYywqpu8YVKIxB7bNFmA54UtAAYJiwWshGiETYj8ymD6ox2JNpIo4hNLE4iAXRqoxDr42L2
T/YsAdTJZ9YUzsT+VcYf33XKOC+WTV7iS3bResgVxdwMhJZTCSXZmYGCKQAynzYIE0kHEJO/ebb5
sx3wIFQR7Mk4WhYwfYrhBUMgeXgtg8oE9RNhGAkHj3EKZSV5d7K2FHARDazcE/mdlDGs+LyV2nmm
Us0YIZ0vGffi/hV6bAMifIAP+X2iesHx8ChxPiFFqoCPgDnK1tGyod/O1UHfg7NVYdry1qRl2JRz
7IRttla/j67W1JyEp+O6iOg8GZFyeb78X+p0Vg6tI8BtG6cCuKr1dOOzvJpIQEmBKtR6dPQzJgQD
Aamh5QmWSF8J5S3R/dBYFVWoWf1hifynR8xVu9zHO5TZNYzx960SnLXsEfduHWNPxV3dtUrDQ7xq
oskMOMNsUHneH2HroqBkGhM1Ye0jkKu4O5jmF5GL8Pw0rB/2TMue5uP7lXjdH2lWeZ18rjOo+dtN
SFW0UMXi4IvDye1+lrUCPcUk4omt1A/wre8jEIxbLvEn6jP0yvVZp3NvFdYMhiXvlOZ+qQOF6U3J
dbIG3tL3YW1MDTR1TkfrAvjYWMaX1TcRUEGldpRLBfCl7dPg4ozQ66uhT6G64FLxrDKj1/sIiSSJ
06rS//sepforX3XM2qiTmYbegesGHpkRUQW46CAzJK8Ba/28hMzXo6SeHuXity5lyOWnwCm9/lm5
N5QMHvEwbzopjBOXLNGZ5GxybCgoQkXRZ/TapclZciedBLBloNBUB4SmCljzZmuVSjtY6Ny0DzM3
rlsuz0GBqOCPeWweUHce6qOVNjUw9Tsy3PVeJr6uMcUBFBq2SbR59pslvp2gqxPq+3+N4HjLJQ2d
Z68TgvXQe9tltSvleA+S0X3tsK+JwKsS7M/bwqg3CinCS20E7KvpImvZ4IAjMRW7hv9a4s3vcBQN
zmLyObR2U8eM1cQlcFdAszG9CpYQpMBRE2cWQOfHyIDEqQFftweQZxvQdC8s5FaIuuVxQyCMRAxs
qcYi8nWsJikzh/jKXGXpOAu6ErcFUu6vZ2DMunx/uysug9Mcj2KFNKpXyuXVSamG3ZreEngdnPDk
s2UxWKjxkuQDPOKraq8sevst/A22k2aFsByk1ZCBE3TEI6yP2xEEE3uaue0ipbbD/m+9PVlMQ8cC
Z69P9QTNeSLoBmhjZszsiWt7VOdsYt/Lx2Az1y2qyW9BtBhAOHIC2MI3kAQVdkQ8laUIxv1dwxXn
HZotvJOIJTfz79WZDCSKLqxaEPGPQBS920d1Ku2mwNlDPpwothgtWbEjEz8r7shML+g68iTPZeNN
Y5kOMwH7stXg/T3wJCFrbRu5kQ60j8L8HuLYhD0keKHMbTbD5Fx9FHi1DzJhI3pqZ+W8Mk6ZSu42
2UfRRPzkvXcwrHUZjyUnUTTtHQ4K4y1e5IOXgYdWqKDO0FuWDmclXup49qwtMekolQPHxrOGHsiL
WSzfDIve3rF8a+RvaqGemVD4tggWJp8e0ipk+ai9CPQA2A5R67tpiUEYzl7/nKcYp9iCEq2AAkvb
qkIXxq+6e2hO0RRDp4c+sYK5z4K8A0Mxh/tr852qPggaQ1wgtRTj9d6MaxcoWWmDGBbi+AvITNiL
pfRdeO8DlWkBHkN+Ie8j92SBnsg5bmnplwzoTWZOWzK03brGSIL2xwyd+X56Fm6FyPSBCOfXGMeE
NqzzEgIi7l7fEUqyHGzV6N1vH+Xi5j7W1EuMa1Ov+iwKrREHUrOp3DnVZ9pbCwwKYAAqruPf20ZB
NhZbxObvXtfeyHVjBF6+3nqPBg5NmyNMlkk5xDXmwtiZdIaxSr5aw2KvprvjvrFAF7pfa7MzoAE7
P7HkkPpLGyFnzn2tSSQXPIq6cdSLOobUZP38+oZgpOn2feEKSkgl5rDguqUGT4SAJ8KTeYNYuZU+
A/DL6E2hBXDE+U13NXdbbUTMdiBK/nDVawgG+/D6gJ87qOQWwXAcGIrTMIim7Up4aN5dFob7AMJ2
IxfmMdrQibnIHxlc5h+SYJaJdIp96Bj+5zlFon25cQ036VC2PCp2SSoAEe4Ywsy6T55ffNFyUo9R
foi00B/Wyps5gCs0+CplkqrBu57E5J5jAH1qZ0oV/WlGNxR0QApTym+IS4kqw/gOrUn4RHojFX4C
Ok2gacuTm7qzo6uzdy3YhfqTzZ4LmM4avA2xhfvNZZjwVE3PGG2yV1wgazF7Uq2945i/GQGZI5na
dtv7xY08PZ3pnjMRsX3U8JdOaN/TwVlzyEnmv8iNXNll73LoNl5j0YVzgVvivNj7aXK0KMwVhvXH
zrHX7dVxhqNWzpQq7zsniYxCxz08y6soTia+Y6nwUYVwecJeCou6uFkeFogmQCh/cRJa3/DWUtqW
0EJqmtGt7+SsME1Flfsw/R6udknP8QzXgnyHLnpsIZlCfLYvweG6xf86b6MAIwl17FKkjWRaHwVz
MwIhzrSTKr6OZE6dA1Q9D0qGNBUQHwXpC6IuUTQcr+eYbnq/khwATH4y3Gz0rzx5Mt7bvptidKff
WYWzAl6CqFPg415H5hUp2mi1dweGfpT59/GX+0eLIj9fKnEAQPk4QYGXsS/cJ/TIHmieDrHc+ixI
ZNPB65iCa4iKhRpxvZtP9sSr/1deTRUreWis52wrBHjI96CU1zlvGUH909DbE67cN0TPgzTR2yQY
UNOE+s7lp+naXK3C8WuGObLR3PqPq87fOH53m4Ro9SIpBQYZ2i2jOpP9hKFZFido4qNTeS/butVR
Pv0K5YPixxs8Dn8cHkwQuvkzzd3CUQfFhe9UfVCJA6Cot2YCvu4cpK2qhatbWL/bn2Noimj2gMGq
42C3RUEzmGdUE+ItGNfHiMBCGSLlcpKp+g4TiIcoMhVnYio86qPX307Cn3KBd5Lp0OORviQRyVZ1
Iy0zO3g+55Eo93GxI/igGBFLRokewrjWbrhKtlpD47aQIWyrpwusazAPmTrSTRQ619CpIUMtYLjL
Za4sxtJwjJ7saleZFQowWNItVVltEMDeaFXlGIPTv1XgRn4Q5mIMTnUdjo+Hja5LuJJ+aZ+aGn/b
CiLrb0vKI3FeLkgAPYlsHdnvdH/cdm/nrg4bp0/UN5h78IHMwQnYypyHGt8sSv3yairvivEJajm2
ODzIFmSa7SdAfDBBW4U0R4A9Uh5zQC7BhhPz6k9tKCeUmFqA3YBIYwOZlc9Wlr6WjnUSM9BSaXXg
2l+TyAMXPLKW65m0XQm9mHkzTMik1OqE6cw5VPY83FmYBj3WB2/OiBap9x9wGbzTPmDQRl+l78D6
VWUqFwIjtMFlW9oJKwZj8XfaIHnq6O7eOiR8xjvpAc7P3QoABdmKy98KvseqLL7IhVPD1bWRFA5g
CXghbM9lFT7X29LlIggsLZDlzpm5Cj6hWqX1ofNfM6TqM9l08oyQq/WdbOpQ10ubeiNnDNcoS7TJ
FHNqyH5VgmCNF532/42joNzyBZmPKwN/GzN5EZd0o9h1Q9YAYJrBBhIHeEaoXitJ0O66G9pGPUf9
MFSD0D6PZsvVLbLlxnodfCLC//qv7HXyQh6YkwN1QQjwYG5WNymI4Hvwjx1mjCiE3ereBwdP9cu+
snafg/URzEYCqp5lPbnVF9Ja7r0Wv/Y7jdPfTmWVMAzvXTC1XXyBEK5iR+2w0+MXLMx0FLBM3Kgn
iZby/dyEos9jQCmmNeKGZXfI+k6Bd2AsLzQKcJgS0ef7NOzh2Y1UFbyEQfw0++dOSzMFegFW9VBn
ZL4I68TjL1BkpNeQCy/lwJICVZBqZWU1iD3HokbxIQ6KfKJeziAyy8f+c1eZjkeSUNUAM/mKXSjn
3uSDBo7YvZQ8FgYZyKaKrO0G2Y2zwySZ2ZXBhyTyWLrxNrkS6kDeEq32raEndtQZGKOBzPg/CM/C
inGY/Eqg//Skmv5qQB+cz9N/2+Cg5tns0fUdCf/PS1qKlgNV4WH+lRnna0mDB9bMa8oUJYvzWqnK
58tEnvtqiVtxRMQpvAQT4U/s9CRZWuRcFdQ1ISv3gQdXATSbqPAK0REGcphWVQUErQCM+Eu7sPqs
8mKKPV4B+0dS+cCiC3zSkAUe1sf2b5ZvrTy3AWlrmTnKYbA7T3nSHpHuUOMvCpLdmb7UI/zPJpKt
q5uTeoxFgYuYGkAFxzCNn95l0mhJdcgE6zJhbqw+HryUNlBu0bxP4iaK0NnR6Do+MFOCKJG3ozz0
HAhnK2SC2w1IW2B/cDXTqDRieXy6M/Q13J/S6iHTDLCJPKMG1KZuAg6G3aDL+OjhImIiua99y0va
9sBjMDfcaK7FMRYJOrgx1IHfMsBkh3qT8N2Vegl9uSyPKA7EO/tFMGj3N9Aq1/QJa3Z5SsxoAWfX
hpwTvofQdr9GSCTyy7GhaHdh1ioh32zL6A0XGLuhRwsoYJChxAoHXUE0jdn6Sh6Fg4K5k0MzirXI
OqgGsi8owG7w2DC+ki3cxOnQHd4Qjodo5jL254I63+qSIhbMIOuwDPM3CS/7zaxfrMyhZnBiNi8B
8kDC7vGdtA7ahH4A0SCQUWxeyrGV4iizAYhHxRcmYkF2xKdXS5yvb3GUbccgoqZRyHWwE5AAv4Zg
CXzJVXAyVYmeco5IVSJ/gHCh0+RG8osnXEbWtEh9DGfGX0vHyTPJ7paIFWy80tc7zQAthXLkDeUb
nem7RH7RH06vh+HZPFzZuzDRIm+KwxYhN4lLb4W+7albprvNdd6S7YWwKiVFUx9lO7hRuvEtTJu0
3XzLo8biBkkixlgW+5fkDzp7LYufBw2JqH0IvJh0xf+PKLkSdDM0sIbfb5zxpajI8cW3SvG1U87/
3FL/U15TSvBFLPSjOfDGgrn7mHaMpcJCcZy8ERezd6n1jvouOfRPpthPxbHEP1Djikjvyi2/Wwtg
lT97SdGAFQhoFFdyBUG7zARlvLmisVVFMAVeC2qmf5VKFTUv7+zudSC6jfiD1mbW58XlsJJ7FSCH
o1QkVyIgnCLEObNawei2Atm52VWPikRuUCZyPJKOkj1u97nf8+KWmb1WFw03+xS1v0senFqwFF0D
nxbUSMD72iy1gJQPXdpmxwJv85BaZ1R7clht+gRJ/8IsRKYrFw03K4EfmqhRzgyk/N42wF5ivJ+r
o1L9aboY+cEAnSm9msWFLZk64iJMxcbcIAhzL+yAJLg1K2d9WdmjNxTzD2QJiPO/i5EesAOBxNHi
pgBvSuMdrjk0MIwN4olfu24W7h+2sdiWhFKky8WF1Znk0jdiVlvhgYzfTSZp1dyFokyN7FjyRlue
1VdXBN1sT2BegqoWxX3/tzqErS5RoYJhG427EJ9cmq/1iu2b7NaWSzd1SXwOvNXSOnYp4PghPhy+
XGq5WPb3x7guTt+yM9Wb4lunwMG9lO9iQKGqt8ZZz2hY31U56goN4z2Cfo5qr0FpdI/sbjP9PQHX
skHP9jbx7s+XRoaSKbcPtvok5Dw/euf2lv9YnehBICEXgJ3+IG2iqi3ErHf9GDSW1zaXOGjMpbQ8
ImcLofMU5Tt6mknI4+CSp6cupoeVH6iBZr/ncjskm5kRkYgSPbgNxZIOhge0vTMV7ros+DJRV0yN
ltBaau/SjGwAG+TTrvF2XME9dKc4Hv2fW36z7lx98I6xTC+2MHypFoOsdOLoyHkRQo8gbzBFoZG9
aMZOCSqM7M4mGTSRT7VBRHx/98BJkl/s6AjuBuZLl+OkuVjpJ4l29NQkqg7pGf65h6qIjeZdK77m
5BYVk3wGf2M4yfkI0qi/6fOH8xZ0+gAS6qbSmYRfVYvMzQhxW/xk2W73z1YRpgnXvBGcSt4QNHPq
szxHey0YawAXS1sdFhV4LhHRhsxm1kScvoFYYoxJtgPy9x2XPWaB9eFvYKY+0zGha7LF3pe8A3B3
+bZH6OH7NfCYa/OeoafydnnoPFkGPqVyhv6MD0jJ0RU0l69i1hCBQPTQX2nRb1czT8Pql/f8xPwc
eCh4aZ3FFjFTe+C0VvP0PXtVkz1IJJQSHQVE0a0Yu6+vKtQJX+82GGVD9BgX0tgCKkW+MCktTgJq
3lDrU7S3JGGbDhcja71yz77xQmiePtUHZGXvIbz7CsKMt9034UM48Am4Ny8411EgRIRRYWrwURcQ
hizmiDVe1mNmgFX5g302hlEBB05bHWnnB2CH6W4kG0naZYXrAAeoqfpgR2IxjoKpoY/ocBX0NN04
4CfnEtaPrXPGD3xv7WlmNIrrEeUESY6Eo5AaZPUPmgcUNbwWoW7JvT6w2ovfU4UC1pfXxArawx7J
e3GOvvE5BJ8SGLswuiBFK9fLnDz4QQwhhTZmY9ZDWYfLwCErbCkI69iCfAOijn3H5kwwRwDo0aPd
76z4T833nwMOAos7valu+1ODGiijVF+NNz96sOfzzhQXkUYWZ5Ny8MSkRqc0DOy1lNuwQeTWOeDO
7OdmzxUNT7viv7nEfWn6C3jevdyJIKaqoOlr4J9SVm5HCXpnGm6bnJMiXhTCKA/BtdFAa5PwV4Bo
MGFWlNYpEjOrqk2vxD4acjDddh8AkJne5u5OHAuClcrcQoFSOIuH5Jw7MnITgR08xMgSCgCuRyPq
/mBtsAY/l7CfPU2mbci1WDIBGUsX4gfaKYDFQVubWc7A9x4mE68oQnEMofreBG7J4Bwfapj5dTy+
Vb6Hzi6qckKn0/bo5I5kAx2sCo3rBbKGSm2Iro6O6o1ktKCYrDFJBpNBxW/5TjwCWeasOcjpS7Fs
zHcyVWTdrNKqn0FrKpsUyjVRasuPYz/e80cyLhvjne6NLcpe2XeBp8qNI9Dvp4sWp1zmjApw1kwj
klHF66oxq4o6o8KY72/pjdQAiNn2Iqd/X1KZurlFYSLzDoPW4HFziThiEmlo7J4lGY8Nm5g8CeYn
GSabpwYFXySu21toPumgGE8XMC8qyTr4+F6DRWYuCCtb8+D0zgajeJjmEa+HWnQiAzVzrHk1hAWX
qG3f6MbwJ6KW0x3XpZEbBTmFnjsRRW1E7LBZYQlqa7hPAwlD/OXDutPjQQuUdTt6Ws8b34LiVjNq
gFZA9S8H/suquhpprie5/oe/6DFI5PrDVYPQQQudF8YNgFFGEFt/AlZrAntKPBKlRS0aX5x8miR2
KkpmZbYcAp2BEMTvLwOdO5PhVzHuy1owxCDb/DtGqXJo0F16Z/+h5oAJZM4j0b0Oi3baVInzhoQv
ZdZtrKmnxgyGRSXV731wnRht9aTfW5KYvqYTy7J5LmYJsEX0Ca9VCbllxx97Z4QDc5jekp2m0apE
ogOCkFSZJzi3xtTQDDUPK86FFX9Y3INccuhCmxv7+uoqrgvTshru6nbLu1EyOU2QJxSRWgk98tZL
NSQcUd7Xm/Fbs38znFnc7e3NeON+YyTXapJ8328J3cz/Yft3ZyXCb2vPJnZ1eS686CsQB7X3PG7y
eqWzGUIjoG8vfZrRtBwv3O7ehquVb8jOTk787F80d6jzTGS9u4zPlo469BTZX/KtTmef2e+r/j1B
KXQet8H5dOfzCRHHG4NQXk1cma93BMyGoXGOPKpUXCRFrRjLXiGpm8skGBkI7Jx4J/+N+wlx6u63
UMpTpMm1JDawTGeCJvJM2C8sxDrYznntwNp9Iae/2wHFMegb/nR/TUlxeMOPSGjBb6ftxqYJ5I9T
soTJebnrtIgkJAXPC6GM3nO/9FhZfsw4i+SJtIDBCcOxlsY7El2w6wq8kULf91EvbimcT7r3Zm0s
VbkSzKP3KUCu0VCP/qn2IRevyDnUKafzJ98GgFgO8Ql2no1bqhgahK0Ptkyz91r5jQCuk/n8yXKq
S77wHIuucgBkklcq7uYesbR2MjyTkqW3aWhzmBtzRDifBa7ySe2/W99t5/KyMe/gzDu9UVfgancJ
HalSlcB+diTTPgaswpyvyPxjZ9K2ck80fN1dWV+2e2/8Zj2Y4VW6nQlyWx3S6YX8Z496ZLZ5EQl4
M89NMitZNLmAQnuZKG89sC21z1FcOJsGJsEZ/LBVEP/fQqwxuPXlw1ifTXAGcytEBLKKB/pFLDLQ
3mW0Nj4sTTfHW7fQv9wqmiSn7DYdBrSKcc1duBuqp0dgO8XczRgijbEPAKkoz7U9jpGZNBiSJFcr
LfiNRdlQVxI0Lc0l9fxRibeJVzxSsJEF2QJJgn6AS0JbarOCY/He835bDPZNS2QWdgn5MPP/iLKZ
WiVJzL5ugCBw0D2IYUKfVjsGHFaNAMwT2WgTb7OU8NtdPgPMIltwzJfP94y4KUfw3tvzeEBySKNS
MXFWF4nLYOJbhv0NvaemTVL5ECIy3uNH8QOX+EFcVUhqRSeZK9rZm06+7w+elf5oUKsxa8uOGd6v
wJTCCWHpwcQ1MNrM95Bt/bV7Hya4Md4iKIor2AwbZKK+hvygCxEs37XcVyYru+5P5CO4AZQKlh3g
42Z6OAAzqgB15/icvaRPkz70mGidnzow2xz17MtlhGiIszpA44Jq/D1NYO3KMlzLe3ZQChxo+yEs
c+zZHdQL6hDOETip83GcHFruZqcdqxsyXGGt005um9Aw9DMxXno7ffJcsUF7iuZySbqpqwxZ0/kv
oxBitQ7Cjn+MIk5V/MyJ8aoLvIx73cCTpzKHoHx3F1v56QN1XzLZKajSh/GzBtXJ+0h21cWDkkQE
q+oMBYjK+s0vVfzA8XtD00j6gswTILsss/0XGjOHNkPtC+Cl6HSU9ClODMLYEJkPrhPwWsZsk89c
god0V8HVRtxrj9RUpAF3iwgY3EZ/p2DXxh6YWtjvLpp6QFmQZ+qkOU6Ow8Xzwv8CkQ5JapKRCoOe
FUme9FIWT7klqwbp+7boWU3w7CWBT9uNq8kjHAlRJ1hXNOBgoP+vc6Km8jzI0CPWlSAL6wWnvvFb
kOJ+AEtOs2KG3BqTToG+2UNbDeFsG/xcR6ja+4BFn4KwQRZ13xTxehiGJamFuhJuFSIslTF9IoQM
s0jAIc0MyYZtF0Wrt9iPftC9usBncTfZikRJiVLrCz0IR1tJtg9vTMxrToV38IZ37q6L7YPsJ6f3
vykVdRHVnEQKLPTwJ8Xt2v2Om7sGGWlsAGvq4yHMHlp1MVn/ZgAIncW4/WGxxYyR6tTYwbWsDqaF
psVN6Se3Fpz2ETOh8MtM1h1X6JyacU+FSer22cQA1cNTw3mr3kEqahTsro4aibJXxGIwZGjwsUj3
AI9zQdCiDVCuM0J6jgPCy5UOPhrHLzp2AMSpXHa5NPMFLj9r4ovAp5DYTjfn9uw2DLLwmo5stA2Q
nqSPE8nYrZTu886h9pOEJ+FCFOieAgbwZRfvwaiFBpSphT9oyZmAbC4BaTIO3mKU1m3xIXaFDP8o
bHf9JK+GV7kHQdPZysd0lcLLkFbzuRkKGqfyiaI9UwwLURXxQzQWevs+ks9KnRJeACwujWghJsby
TvIJ0fg36x3OGVPWkO/1py7Gb8SJOPcUlh2RfZ7OkPFYOzkV3AJf+mm8sflSr82l5C7M3G0BbULj
49ypL6sd51TUSoAVlHY8sTMRyI6TKsm0PDI3ikufG/W7TXESYJl/1ZB1w+i7DZ/8YPmDr8uXXqlQ
PVtqJUF6fqjTGpqPRKjSRXyO/B41bDkd5fIAHPxaamOiLah5oXOAjTMBY+fijMypzXfDijKTJnbz
mtCoo9jbrzUNkBfhFLmAWPOqzRTpy+yLCL2nRN3S6e6a6hdiPan+rQdaPJZuUR682U5plQIjGWtI
RH101ZvqgyN/NFyjEMtqP2V7sSSxO1Ob5dSO7EkTft6M3yB/qdiYfy5CDM7gyXJBGjIjOanLM21n
QuNT2WpR2XXHQryOJJdNUl+0Oc4bzMC4yyWMrGWW7mM3i8jnWEC8hCwqjxpZxto1ty73V3Gi4CaU
dKpsrGqR8VqZsVeyB2P93woB1UoSj2dNZXm7NNR0cwagVvVX9ZiwWVhKYfuHutcRoIisZqt5UMuk
4ljzQTY0Vc0uEUwxr0Xlwi9Ebo8YMM2LNN+DPt2IrTotYwGwap2UO/ijYD3zIDhDv42ouhcBesyv
r6Z8hiGADacdcZ8mYavKcEOIFNppp0bAMHDdXeDdaPRbTA3VmN1Ky9OpZVTzlBWgWeVjVqu0m4GQ
z5cwpJ4sEtB7p04gYFNvnqz6K9pDNdGbw/4qO1ZptLs7Ha/ZdeDAX6u3YXanFXMWATklWtxlSZmF
5S602awpfsR+n2UjhO+hmIwiWg7xjuKUk6PhXJaguPkzzLMBEtO82e3w/OHEzyLeswZdDrP5UyxG
uNMixAH3iQaidWTN+ETb15A17WdJQ1yJLQGOcuxHzuO/TKKnqPmkeonocjv1//WJX0sKunz5VlTF
oj9vsvccLZbkIYHdhf6rLYmGsT1oggaCDYM68aT4ulLZkUFIfN6VWdvYCj8T3oIoaOtvFAbGcPO2
CA3e4qXGPl6+f9kXD1NpFVDgLCuYCiUzhbQRFQY9lppXTqf5tz6DXiOb1xAm/+/3igLc3t+6+PPt
e4kT8N5VNbJveETzQ/jSYjUMLr7ZVqfkkAJ9PHNF5BmWBEdbuwoVmTEd4zhvcaof+dQ/xeFRW41j
Zz9xZYA1gYq0NKQT4LBbpkMySxxe/C+WYj3eyHp9C/spNRVkeieVZtsJFU3MdWsZPVUekPj+03T2
L93usqk9aAlviA8+CilxuhGWUhFz1s6qhVYM+26Mu5YpbXjN0dkrPZqOejXlJauyIkJmT4NSE8qT
m251n9YYeWd31SMx7NDRxB6xUmC+tpxbHe4i9/6fStuTsWwn9YYd7c2gE6XrZN4R3pj6JWqTX9PP
eAtslGntnzgzppNRwG4YWU1o1Y/4IzNrlYFOmKjR9eAiZAhb+s11ei3lYdzuLOS9TJszrm6dbCaB
fI1Ca9xi5GCRXxo/XKfXBNz4fNOy77ANBisG+SckIqBPW/ENa1cN9vqPApbBfzTiNS1VCL6KxrPT
3Q5Cv+xqWY0oSfCgc+bhEFtbz8+krslChjFwBj+401UkSR4gDBAehqpSk+jFVs0sMVeVHwSA0Bd2
QtrI0vclZ7a16/Ar2zJT2YZqZlffjs/dkqOPEx5wbZhd+rhpFjF7SUdnwbokgOerO8C1eYWOM1ua
30cDg37Dh8wHo9gw/1i7nSjAheuQGLkhNoYzThtyZ6Zgex/2zgCqcnAXlKB+gZHGADv8lM9mtEa+
YUz0+40wJ+iul/zQNC9bPn/alc6sgzUJhETfKfDe+sShk+X/I/LDEmywCD1byBcZ3TI4ww2Z5Jqx
jGhyee9ojQv9+ge3F+pWpV4eE5DN0zuPyNLA5NzzifV+LpH7f8kC36vdsaqbf9FW/f6F4NfDIMb/
xDJZ+d9mnTNiasCpBpiAngf2pY7XWCCLzixkp3gwEHheZOpkrpD+/MDOAnwN5zrE2SWVojnEukCE
1KtaXd/yK4D9sDJyIo3yrkV9rBG9DPU+ThuccypVSTVEmfXbHVwfrMkq9t0idvv5UGn8TnYplJ5H
/aXbKhxaKZlyt6/g7jOEbIkpr/IsQwfUItghhhRhOxS1LwuQe9G8z4NkjnMZVqmDCfKJHGISI4SD
5aAFFiWxxnbHtNkicVbNB3fahVUXjOEHNGUyjNJ+DiagMnj3Fqg1R6VGAOPtfsum4LrF64WE2PUu
tuYYFVmqLm+7hOK7JS5OuhZGqjGft26o+4X83Xf1SwAIYLvOrUmigDIJ3s6AGsxDarJ/F+Obq7vZ
oBNXL/Rd3e169LOEK/+XCMs7doxvza/e5x2tKolUyyn/n2JtXjpONeA+RiePwXBxiv77P0UGUV6j
Evj/nwVgIiEfjkdVgPGmQyfIlGeGKul0kM9Jnh1S4taGyeaxfJCPNoX1kZxueTpc6vZlEx3MP9XA
2LUMzbO3jeSZDcauNIBES0Om5IRlpcNlUuY8ze/GjR9sTKbtVVyyFi22wuWdt45ol7j40RRTrqSQ
20Riyx+A9RwNltZSH9hQpWjKa0Vur3Q9VAFubNGkCxnF1qshHKjbdwPzi3m8tOPDgdnau/1ZVMkh
niProzU7MAsjAcTZNDwbGr2LZ+acANn5ryWfOi4WDjF/HDdZDbNO9Ob5xR+G39HTn1J9WodfUFjp
6Qa6GMNg2FXkMCcZModPE44Wl+cKQe85QeyeN4lOKovweoj9vH2bwblzLADigi71qM7E3+uAbRdH
0bA/y24SMAv1pZ1O4WmZEgXTFnJ4qU+f+NyKnY686lBqUbYADAuETY8q1cd87tgnwOhVuj52fKf0
PHbJgKCA7JZ96mBlzUQnou50gtBidBNxe3wsV+KbSPsr07f3nYELWVaJmPJVNdsZfjr/Qh34Vpby
sVZZJt7Wj2cGBW+6cpGMQ4xWRWKdb0qp+FO2CqmG0Z0B180RVHGfpWJ1nKjOH9lTu48Ok1EtoqC8
sn5XOx54WtHlVoxOYxKd6JFefRR83ZlYRlJqKTGe949FzILUSOvi5q0HDIWQh2+arORjB8jfEbrc
+wUQzlpZCI4hxDchT654XqDe2mVLWC2JjdgO8sxGEOyTshihZip9jxtZItDLC5F+30ntWGlXboK3
CnI3rjKe06sJqSE3g6swtFJ+0TM9KAWldLZohvz3BiE7FRG2ts7tb1PJVr3lL8bm8SitZeV7Zz4L
KzyxrLASQ/XuUM6To+TdFi10g5GHxDcaBXVkIcfvuK2qt/r2I91SYclMdeZBsyhsarEEF5oy1lR7
ey065K6LPzr3EXCb7aCkyllVlh8f5b9k1tMyCMljI0r2utZrFQig6VLWtzWSy1Neh+Yho1FhT4ju
+6A8q5Pwt9jmxTW2XUUQLOH2Ihk6GOElupHnL0fbwkoFyrXaI2y4fxjCcta4i8rW5YbMGInWCrPp
s8Du1Iel5CQhqHZv4mxLCHZgK8fFuj2ldIXshEbdQUmdccOECaVDNzE/JRNUYcmB6denfmg0Q0UD
T4BNyjTPjBbhncwBPilgoo0F/Ayy6DXa6IlZPzXcC5PJqoAsFcgt65NWJ1gok1nB5ju3eD2vefd7
bN7H60oFGt2IR/Yg2rAsr492fwNWSvu+oBKzQ9fl5mg2lu2LjPqXne0QZRhJ92g3YZfacg1RvNXl
9uwn5FMdM6I0/ugnL2Yg9QuweqFSw5gHk6YMlnQuyOxxU9WGBqaCH8AZdGx/YDFAFaqinx7Yxinl
bv4Mgq/hXKG80liRgS00dngbFDYwFkFi02WwuOd6tlma4R9uyQ0ZBm779j4fy2pu7+5Gw/f4MBP3
l1cQvjsj9NdwfECp+94h8dyUGGjcehwfAHcpo3aWbtdmg/XvsXmwgM+p06SkRxvDQH+vsJBcQbY8
L4PtWd24E9VK8U8d0EhnhNBtRMn9fpNoay51xKpFtgsuGww/51ROEdOrD9HB5NV1j2nztWuhEF8F
KqjvkeRg1qh2s7Ws1zUkYL3NnnY9zpWRvKj2nJ7FlZfJNJS4rqeV5fzl/P3XfyY21hseWhOhtd9F
oK8Yfc7KeWMnm0WY62D7Qa3YiB1Fnp/x3Sqz8Eaf595g/x7jFscX4RXYmDkQbOQZELbvR/RZKh6T
Yu/dEyJTsQIkx/vcNWiGxKZLCioOXgv7zMKIoN635VLVTCPPLUrjkFeD6huXRKJAIXG35/BiaCka
yoYXRsXiMxZ2JOcyPHPLa0QC/uDMve/wDALa6Rs0dB7NjvxjdB4BnJ8ftAh868uz4YiC293XlpJm
xtZPAjO6uAa1KUjMXoaYonjy20YD2AAAux/cIss2cPNB/wucFtXE3KJ+hgbBE9NLzFUlKwq1Aiyr
hpkY2Cdc5zTx64XSpAb+8spCibbkPxWNF9dLiGsD7TlOIF1Fw5GNECnMxP1TuFyed1kNz3N/eQE9
E5wsT2XGqr8xIwOHUGPONSn6xjZ2cOJfN4Q1jqW9ZU8LMT2W6M83YUQfL2CsaDwBJ1g4uOVLWsI3
ed2RQ7MrFcg3H4j7VnyCHZHrrkaYbKAPCWKKhvn+wzddwIE+om2SWUcUuTMnpUXffvGEitJ7Ne8q
In9hD6r97brInKJfjG1lteLMPzi6xECvqXDydfnLSR4TrrS67tH9waHs1i+0EXuoURmRlOSxBI4k
fuA0b9pCHEzqbKLD7Fjexu8I9L/rco1RXa53cL9gaQ76owv/uV9FLtE5TWXywDabUoG2UiNLzMP6
08Wk6faPmZQhl8NGjbnWxSQbVLdA25+5nmI74GOv1vY30YVVe6k3iH5G6QnAJrpDHGUxvu1OpTZ7
vwqcjvVyNPR92cJnAaypUHFOfHghUxiebN7oUrP1vC6PdpG2zqfhJggXf6zqJCPtXl0twBgb4XvH
jBVM5TJ0nPDAzHcGOJl4NoZONmQ+8dGbNPiA3GD9FQQmXyBJWYtbAVqbxu6PvDDIszcPO2oGfYUD
WkgIKRAtEQ2O1vXg7VScRa2K5HLr9vhk2dXE9LHkVT0LOTeOL2OihIanZc1iqXC9+ocCIHp+oZGI
4XRErnBzSnVIJEQEemslT7sRo3H3MBpxboIvrAtlAyjVBwefI0k8zNJxSNnNIk6mVzgqlr2Z/5yp
twjtQtVsNoSYXrK+uJTFg1INVhBL9sa5Cpmvnv5WadBKqE90c1y9aMPgCjfC4TPUK1fkSl3g91Kq
kCuGHw6A6dLv6s4JMnNM+Yt2YcstAFL4kTjAwOLbxcnFniETHQ4V5xcLP7yTtWSSKxIS81lkVIaS
QJobchbXJgQiizZlaTkq3FNppo81mqIeBK0jbSSs8wdFiBsEfTEusIpJViPGHyObBEC/HYyPW4GL
af7/QB6xzFepTTjtHgT489ejAdQxbKFk3o7BlfARPNg5KUAHozHNf+16llS7l0BR2pIRGYVJXn22
4swn6aWOp5ZtxxjnUFKMH0rjx/arah3GTwtGAbYIOIbKYcD3XZjjM9ZARIeBkPfnKQOb1EWTgq7p
+c1Cck2XZ7WNhip94ULty38TQuLIpParbn0vbsQ/ZdJM2lxEfK2tc1FFpbeLyWASALwqzd6aP13Q
jwCCB/KCoabnXmEyLCWCLKcrKurjLJL7jR5ZrKprXr8YGqemChZHiZco/mNmLinkZizgohr/FjQU
9TtopJGF0zEnSb7hl1Nix1tv+KgLJYi3a+n13cL9cFon8u+YMOaygYWTuWnl+SZePnRjLxAZvaVM
HcYXLD+EWlMZqh9WIa8U0lt3xaBElwjz5qhNm3iGbOjbA0X9RZzmsTxL8pA34v/CNh/Z1ZnAv9oh
Yu6rloUteBbReVJ2oTSVCVNTI6yhbXQS8S6txDJAJiqdyV95udekQSTflytiFedTHxUdESsDHPOH
69YqpZSc5oycM/TUffctCktDZdbqamxHJfgCPY9VsOqVaTsj81aJAWCbm1mHfgnBsRlmuPektWBC
ICN7VpkM6REkW4gBlpRidMR5aOvbeFQeD2VCfzKitP9yKvtGWJo3B4OH1IOA7CUIxt4m1aGzbyF0
j/djatXZAoIavPYrlU0q053eWxeIcgT3PCYHvblEoD078yhjtnknsIQ2/KKykVe3OBTop8j+Hm9a
GYK+I8q96anGGOcZn0PmA7YOrQJN/ccPQzKafBKn1hhohLhw6xqOe1J193tP2+wHOO8KBRS8L8fu
QVocIFUK7WV40lLCQU2AagSvM4/P/VslUPltkHHigXa3xR51UAjjgY4/K5RaXxsGBdZiZPjQDwW1
IQUOx1HqDlFLQ8042zMelDhgAjg4NLs3J2WhMDgRfHWEDoZHs1e91N683YdJjf8V+WbzQRBwQ+wm
j6ujjbN4De4dkP+kY8+TD08zUim9ngccOSO0CDRFKpjH+1h1PEVaJMUN+Uy1XaJeL/rha9F9to3E
FrcpDNnIDOeKLBdqK/vamboaTt6cKE63YUV0ETITBICXHoKjo/FC5ze+wyLAw8NGMgZ/a0mOPkR9
ngzllrUqeKWl5i4cNrODd8g/kikEcDfwgSjT9F1rVwu1Xj8yNKyNb4fdHFIn+tULPBq9hks1C/8b
OawnRjGc7J3lRYyadkAD2Zs/RvfgW38fpUvqyMbJKk9njjnZvX7AOIzFd24AO/AiUq9rDq57LPGF
JOkGtX7hSZER0x8N+wCF95WarsFyhaHH3fCDHdcAYJE5/O2dI2dCbfAv5amvk6I21tYcAEr/e47V
X1BZviXLK5R3dwRV2vOVhp4K00h/k3ndiWU5syVV7Fefis5V53k6JFVj2lxACcD+/gPntIozbrvk
6oVtYiETHiZx4TUh5Yeoi/LNeLPVNq6wXa/F0ra+VkMKg6BtKQhQuSr6FGyjdl2n+i+0YaBbfJUh
gHnX+E78Z3Jsox861X10bzvBqgVX/KCC0ZJakrVH0YElM5umuJnz/S30zYXPHt4zkss71s4Ftgxr
pWIKUtq3Q6GM7ixNse9MRxYsrSS7NMICSpK6HXnK2/FCRxSy9Kuk9a5aUBuE67D8rrLQPu4+FzkE
9SwBe2WX5fxlBsBGIWG+L/eIXS8+SI10suJ21urqMzmSEoijwajnxXNJ75IsTz24+JZUdwi0tdIj
+r+7iKpyEswva7VUfcANE1QV67NCHFjoBMnaXtWHlukT3mymp52eJ8tdfRQ0/z37Pu1H0ob9fckm
ByDxcAJtPVQdTn9lgkaw5mB4PKREdxygbcnGHhrWr1jPq/QnTKKRfX6JKzJe/5i/WbWrpsOk4E6R
vJ/K4SLoCkiDNTL0KAwZsdi2ZW3U7z3Y35OaK+cSq2igF/4FlUMZeaEXsDmdOCJQILeiZuvIdPZV
Y7mR9lBtnBcfAnXc7sK0Tob9jDOdzf2XgkiwHlkXUVLQUd0C9LkQqUbJQx7V5FOMR6sMutniKX+y
ikbv1CstM6Fjltb1SVIyIqep032QbiYKQI6/dKxfS+02FIcJoSgPxjej0WGP31ahj1y4UfRcS3t2
GUGRm0OmB/PHwRK4hkajaTGv1/dJdWGFTHpLL10Y50pEOG+s7pObuLOalSZYAPMdeLgJHiG0dkIX
jULxVtcm6eP/DGH8OMWpK3pYb2vmkJQfhkyLDplKYY45BP0qBtebZk7G1+gxuzi9tojaQ+FFFubx
4/K4kyXKNv/aZbxEgmSmOJuisiU6EdT7WeLINrdYc9ADebUqIQv2mvLx7T5V9M2n1hBEZro1iI8q
WRI4ebGzJznQFuRf9eBhbiJWypBQYhgxi6SmkvTaeIbcZL8tXA5EJ5F/L9DQ3h09Ed6dRXVurDAo
xVsKikTJX3vGYq5Z/Jq+QAxKH+JQx5DEQ0lF2yOiJa7d2s1jOoazDBfA5Z9ReWodRgbxqUL5A5I7
b1KKZN0rfUT5GYSPTNaxaQjxrJE4oCf72nxyVYtObmKapjyx4zPkaUR8RLokAL6S+it+qsxutWpW
2PPB7sG+cUGKPShARBYH62zBAmFwi2clX/ddRx9K23jVOdpXpk1bMpUGsfNyy71vbd8QqPmwJBVp
i6gTZgLjC7GDZ8GoBgIAMUB0NgQl7wcPaxspbnUinRXIE5Ntuhg29iVoOrqTQQeEs8K9eBw3EXZD
Zv7uiuwsokry3RoSAD/vp1ajw3BAMqONGx2DH5Um3VOYI15jO59+ICe6nWl7HL0nZUYeognE/jKq
JPlCKnD/9GL4sBrXUXSH6fk+XKpee+J8pHF8jXm3MU9BoJ0QJupa6+BHxaAoBNBIvW5Nu9fBONj6
+cyPhX7ZgdygfPsjrTxZ07UBXb4M/anRGUlDkTnQ+oSLxdsHedGToT3jt1a3Uf29l5ufWWGY5UG+
6DchLowi6+r1D26xrK066AbHDxegDE+zX+JDYXYMMR6UWW8fpaSAxyYM88mA38NWmajJDIf+aKQE
MX92fpGkbnyC1UQDhfKBQtQv1Gx7Olt8xVF5j1oSq9Y+GSpYB+ldDg0iCT868sRuvX1xG4O32Jln
dpn7Tt7Tvz96tSFtCAQY4rNvjQAthUfRf29fUvO4zvJSObMDD8zD7B4cjPi9TQ9/ikaagSz2b6Ma
L57LdkGB+q/0tFZn6lbG+vR1ERfdpbtNjHYN9juxF/7pTGuvsyt54SzKdubWzaJMpDe5QbCDGJJu
5Z+8mg1w8yE+1vcUxPGzcqCWUODV1hKZJCPP9VNsRMYulmdSvkDi4/QrA6dv1so3fvbJzt/WxuIR
wmSpzoDBEnwzFSzJuppfRjmyBXPC2siD0SY3bTmD7f9YpJ2E5Zsvlpqmem/rmNLKwnN270ZSTLOa
AzS7pwaGwjMvuNh5zT37Zb+qQt8cchZMsPF2bOdotNPexQs10M2wK0qMr44VlfUnXLnd/LEzVUdR
AoPmyUKkQ63xX4WlJKrPW9XiNU0xAkmGYKK+rhgl4N07ocbUBoh8GoyYJLWpvk67DQkni8jgaucA
fjZOppgZXXr4stkH7HW8tn+ZpzkjsKHGISYo99ZVwIJQs6oW1pDPXEvLuQMP36mONo45HDSHTvDX
aDcAla70YwqvPZ2cbwvUWWdlAHc6ssr2q9q0CkQ0vJ1/vOUHFg185xJA0WrYd7FA5C85KkvqfblI
oi+8PuGsZhxMQ/UujbsyXnBygJG5FgoYQIe6KtPP0Ds4Davm7giSWJvoF8VcjER2zrAghtvlp8sn
Fl+pQvPUqn7BjkHR5LDdGlM4Wr1wWnXYnbrlcHYB/b2PVFfTSM22XMFwxGy/IDfrRirq2VsAar3C
m4QxxtCfHWsl8kmTpBsDOpsM5KEKEUNL5uvTqBm1ddBzLwK7tOfmemiBxjk+bqteKQsv3z+gW+gw
Dyqok4+cI2lsJrxRh4WxHpJ2vG/K2859588Lgfa/9mHJlnsoVBlMUxl6J01Jsj5hKD9pYpV2jBYp
87b7iEbUKhEtYjf/gUBif8kKYaIb+yrGw4cznJKvephtPwyUxTshbpVvcShoqbTkVe9zxIqHzTqM
9H+NYJkMFCg26OcoXnosnpd+kbvLnUJH9RljLkI0K+XI4T7xCa3yzowuFcE/JfdKy+VNcAtAap1d
ecB/+HJd6BF7kLrMNx81VZszCKuLMOlHO+eCrTgODmaG83T3H0TLWmnGkrikPsoHzCxJpBjs/Lae
q7cCpLO9lgFgAgFL25To4b0E7vyP87cwqh1czDUxxdsI+PAmcVgdaCST9lDXaKDGcisHSyca7OIA
2rzyZKA+bwP17upclkIiMzIECySKaLt/AkVkFUMiYDRQf5dSn6YKbMcVU2ATkU0+TQPi2747kjTy
8l0oXH4bQgTloU6OwDqBnBgz1I0divgsKvCcuLGEVrlaAXn9Nobn6WClzJw8riEE9mUsUC9qYyLB
3JjqYWDZf2PsHlSDYGcje2MEuA5/ceKIMBtjB/J9MremzW2MaTxIM6AtwLnJap+nWIk1Aldp87Zs
2WkRYW6tUz5okgOJBohQFyTPUHFJBHTWdmYzjlIzsuA3VK1w6Y5RxJ3DZjnVpvCi9X7bSE6vOrtI
BjoVOgj0T/WVMPaEI3GH17BDSiB2CGSiz9wBkv/c6RcHPRE7EltB9xZpcoMUp/KwTMGGhSSce6YQ
KAppmL9zp0G8McD5lBjSJH/vdQXfK/nS2DhxCgmP76w7VNroKyFU3sBHJueumMPIG96Rem/sz8EJ
SdS2MnX/ROK0Nfy+pwvdT4RXXjORR94VEGJFPX9ygd6woa8dNctG3/5KD9JDAWORhRDJx11H9lhW
BqrAsewbRbZLGtkqwecddqPdAZ8nBUqtVCkkX/OSp4tsfyKIExFOIcZgkKuSSwuN+nTCjJlXgmeA
GcqAWXReMvXlFFIiV1XfJwI71DCt965329/GJ4HVvvcx7Jq3z7G4PyP3EwG07C7z2T3dYebvZbiB
bpbIxGZtBDekJoCRw9qPr+kURj0JlWQvbcFftJIkIp5eiVVbSyrCjEbV/dCyNP5u4F+I+wiLwCgo
t/WTEteFia8vazZscs1ZsB6pM2/cwJ3bbPOud1aUp3ZsY3IQUWarv6Q3ZDnay/kKcY+Brh2C4Km4
06775APyhIfUCS85nTMp+2B4Yb/jazVUe1ZKxzMoFZLmi8ZHyuzVpKfoshJr8fdtXXFxngYrzy0P
WUOomfdWUpbyfFdHNahZER3a0l/Z+ICh0Z3c5W4rfGTnaN2V7Zaj6AyfbEVecf7UbU3DG1OY+5mg
Psh0Uese+QjOHxvNhNbvIvch/oXKIPy838TIA5cL8W9ytohEATPwTzDLrc4VTuSr34ZeGG2VmHfS
vE5wrcN9f9f3JplwPrnu+gmeS0LKZWAM9m1A56oeIJn7B4mHw8ZQiqPi8xh6NYWgqoU8q1KsCout
vHklu55kJEgovZpy2d5vpsqHzSFPtbZ2wcPS7Lbl/p0PlExhkMTfEnMoSi8iC/wiJsp58smm+8HV
p80ZLoNa9/uLx8v3JM0e9YRwIddsORaucriBathPcwggfO/8qF5C8TKJ6R2zrWV584Awy/uDhnvw
787WD1qpwMNDKrx/QnxEtCDGIyuTDKGE2+u6tQmswbQkAjTHMioa5BcgfQwkQKMZuNfaVV0KqqOd
Rzq4pTmfdeCbUGwzGev7h7Crphg7042nPbPKLmcc5f9PXmZLVI5KjaEiFQScNUPx6TRDUFGHeYoQ
QNUnmDqs2GEveBxxs9u2QN1LytaIabcHePapkgLql5hnkdxvJlDZi8Koj4z1+2ocNyqfck0hsd34
/PV4IImZE5SWoUow42gF2WnJLB2jItvKBukJYcyzt1ndz8bmqzNjR7eW3qcbxf7j/uEXBbztY61y
xtFGhJtEA8dXb1gqd2inJu7NuxxOVm2afXjPxFrkt/0lgEvONliRo8rk74xGQrdo1KiNIVFfRe0A
G6Xff2ZfkMzkLcwFE4QvnTbYK1NsqS3wTe4J/nvNU2RBfchzSTA94T6pgZgPF+8WNqZcgG6U3Ef7
dPjLI1JaSINaP4cBmVtu8zXHEpaOqcUxinlTnTETr24PMGLRdp+YPw6JQ+rkpU3JgIsPeae3/Ok6
SGkpBGQTAURq4ldiC3UlzkAUec2NKddUVBP1mrOIY2gtN69zYiNILSzAWT7mOUVEEIzV3Ch4BxrJ
U1izcmHaaiC6lBauV632qQJy+lK6K/Jin5HtEImLCn2j7Bg5evNuOv1pzqp5JCNHQmzMZomqcQCV
UUGH63BgIRRUQS/YNmRihTIsn65pUU0KmLBkiHC8gRGnSVp4Hk1ERDakar+bL3gGOtcnZryzXSao
8CgGwI71KlcjKG1OVyyh4vuTk1TzqbJGMw3PQF+8Pnl01mXDUNLZeWg6D28GHdD2wr+Tp/21S4JI
xh/NWfUlpkpIgC8UXRyIfueBrQhvuyCQVpIJ3LIg/FPfp8ENTzP6EbTvqKNFIKTgxC2SEUVzXcQp
W31aWoLcek9ifJpMIgfZIdlwzudWR9e4XDTv5Qk2NVMqfhHRUONaK8SL9aN+IUhg2OEi4WbFip+B
4JctAI7sBmht8aMmmkHjaGGm5vqAz1/L6OGmwuyW3CO0lEHawT9Q4BKcS7axqz9cAzWsy0wkL3mc
RJDTJYrJfD2H9G+ZEisPJ72Ug6xNG5J7UsCEloOPuLE3JktAuWkatVazTZnU6cR0kc6bBBwxmrjq
LaFgbXfndotITOtn8Sc4bQMYeneaS0sLEgmF31WrayQh7K+N4NguI4c79wWRja4+c1/MKCsXaBJF
iM31VaGdVWV1RYlydh+jPG5PJ4nr9rWhNLLm/SbJSmbZrFHY+U2mLLgVW9GVHAsdgeZjgmFZ8q7i
vIZeXsDqWbqurRcWxn1qjOAkxAlbW8Z+lJXKV6FER6/oqodo4uWgmIqjJ4LJ7iGJUmVVTSmTRKrd
AxYRkFM3V4IwKXxtN/UVsr4AzCbOfRIrgJkRIeGBeweSkjqccO1DxXuMofdeZwgxeHA+88+tBFJ5
rxAjAayC9YB5pPtxX/s6CGgKWEtCH8ogtFQBf+TL3ufuX2LvYQoi/FypA22DJ5lb8TN2bHp0A0G1
DWLcxHpGCFpRNuT4tIvgi1bdqdZbw/wdvNGrnoG1pSSbeExoEFxVdP+DMEYR1EfVx3Qf9ia4wNEI
QuYtYJFlRPc4gyyhMl0VXqtDHmAXcBJPncOGQPegAmggb8em99plTniQHVpvxsm7MyW8QeMoGqrn
kmJ4M314h7NsK/WO3wIBKCaY+hnxd1wv3bUpBanRmqvFKyDFKG6sDKmrd3kocg/KyuRy6pp6mTiK
vsAGuhKC5mHmTTPQk/B2ZaZN+pYGEjlOI0/HMbw1rIVg6ylb+ZDQG0eQ5ZGMS9mV44pUSMO01GO0
aarqz75whWqERtmH30lV+n+0qXl2tcpSakCR9HIpLXhOJ2ynjABVnNeJPqjZAxahMm5iEOqnIy7x
NiasLUkSEiFGQBPsFLfpgYhBVpdiFjnG8bGIj3jYGNMfADg5kORmFE4sq/7IZVFM993C1tI38tR0
QrcUHoARghpAPQ6sT+/S/9QMLpCXyxMBScGyd+9xOVU1HOZDimTdNZ9uB7U2s/aXzXl4EHBoPF7Q
n1newEoD6cdxzlZyAYXbjdNapSwF28Yn7npLCLDfr85Vzirq1CiUo8iu6jy3ddZj4Rz0PQvTtorT
qi3Eau1t35iUwjWB+jL2JcVYf30m4njB086izLNZPpR8xlRnfsTNcKd9SMtczFrZeTPMmQNJTeBL
tG+wKRZWR8DMoiQm+R5D4JMTM64pPLssd0D5MjBqvYQKBSMxbZUdXIkHRv07QKiPu16n7pX2Bz6f
HSsYQ8bZ6VhgtU+Gz0adl8xpFdFQhnuQ9+2EHUSultDCx0zxVkRBgROLGArJRAczYju/U51+yDKN
PROutjjCyMsRFDDweUIR6Mn5XmjEIcbWS4N4bhSBDqcFlG8NSJm9UvTjsWxcBY0r3RiASLIAMESb
/xtcZnLuknK4ks+7RYwhNzpjAZIfC3xdnshANQ8SdvUCYzPB2GtVIY1K/zU7/+zyi0fB1YoQvclL
SPUv/SVoFD0HZpRIuU59wMojn4DCs2rwDcy2VVhEru+YiM2aVxFuBs+awwEAFBbdELwtymlsMOcF
zkL1C3NVAsjUeXO4YkkxBWS8XERsx1tOFMymm1QszA9svOpR6bcWL1Fj7Pma/8PjgDLmQ7JIryhu
gtSI7/A2l2111N1D82RYX/txW7sQlUnzc3+z9U93mK27UHBjjwCig+93ymLtkj3B+t4o1isqvRU3
5WI60VswI5cIEEnpTvs/DHZGue863PFmLxG1+hBXOcDatXXAO9WG0jyq4vQmACrB/I0epg+RhjtP
98PzsAB+OyUjWYKpl2X2RkTi7vqiwPbY0woUMWaMI5obFdki0K0moYOa7isaHsfSMXjAIns7eaKC
ivKGrwG9ezgy027TG5qerzbc5NPk7+9t058NPQ3Qs+FVJFTIDNmRgOgzDakc99yUNon2F7+iw+Ly
x+lFdXM59vFgZrrayxvNsjevvOWquXnmzZET08NDK7iF78ErTvDmj7F4twBgIsvfdh21lhqs+KDk
BZRXgsLGnHy6v/Xy8BgKgKdWr5oA159YGY3g79MbHFc1VmdzbHVBQTqH/ydg61is38VQQJXRyTB2
y07jA6Fc+0hVCZqv8kqvcjRFAv0jmRU0MUQZkSXxyKMdAPm7H0C9773zNSJeqSwBXA3QQAO/wX+A
7GS+NsKQv8pEvSCFC3XRBnELyosuZk1teHxuvjNuLkQqb2IVOJq7K7mHU4hKwr+9Z9MKFTEGWav4
7I9ElN+invjjsBumkB7kvDvxJ4NytHL/0LtGJZs88wxlQPTE8/uondy+O0ZCzMapI3ShiVI5mPD0
qWGEq8yZge4cxeKswCWSwtWIzFCiB/MAgOlceeeotfT++GGINnTy54WTbgf6+WB9W96eWviQQRM0
techM9o0W6Mdtvazj1212zEZ+ISIWvuDwTE8i7rlXgB+LSJlEuyRlovBf+WvJr0FqGh7nHUj61ez
1X5dAHiWJ9e2KTorH1w9gqLVVne7hGVhSDClPZssJX3KoXxlZ/spZGoBtRHi/K8SOyM3+hsJbh8s
fwcxl9ywccJt2qAJphLQommwUAkFacJ9/REeKHKyy68x6j7HNqgXzukYfioLDREqvYLJci/7D9oG
2cNQN2hF9zAsAaIs3rRtRegQrRh4hsW9Cd4gcW1Vg6rx1L4Qov9YmTh5rmkN9lQbUznIIPog6faL
luX5bptP434REOO5tlPsDcg1Z6ErPpzJo7xmsXf2Onj448rKrq8by5ORsZCFF2DCQvHj8SMciEZ/
ThlFLv6cWTygL71C9fz1j4jDUMkZPgVV9fFP7tbzxAgn+eY/rtJirm84JtuINvfW75WSe6t2ttgT
QmODMgPziSSHXy9VhMeVPNbFUYruK4Giq+/gcYksP78VROAu8S9E9XzRuMt5JwvZKJaZQ/7i66k3
J2q4eDaflTWp/CvpL4wbxqaxd0tr06J2/+LkM+EPhglCHhWlktICHZ+ryaRWZjuGGvzJ7pOqvGsC
aQxm63gWmS0Eq0xyLjdoDiUuIA4q7EmBGhchcXJ0wiNvu0T0KXBtOVwT+6r6QnwG1dykXaPhdevt
uH5+K08aJYWfubifJo4ghH8ISjBgnO/+/rNLG19PteLbe9j7Z8TrBfUygVeiSxTYu8KGS5xzpqg0
HL/P9bUHJhJbRCA2xDP5eE/+nW88XXxm4tva6AWhjbWnQBQqOzkeiGP8gUb+ZpoIvhOM0fmnBAWx
wZaN+Hgr8hSq8vPeKF1KPzX10j0bKGr18URJ4GYhJnpmb5VTNycd/YNQUqmJAYqXRrI6avfnQCvG
+lPBvj0BBdqQgtqAj+Iy7GBDh14fdfAzua+G9fhUjNPROdNiPPEvML5qu8Cq3oHH/7j1EsS7uGK0
upDbNrxjMRteIRKDqXAArFKzxWkPEbv1axYydDOHU9dBhMvHrES47cxeTLn6fbTcfZ/y+AWPrjc9
3+WuB7ZnoMPhMASF1aqm2NPDeaywh5SluankE5Pd/joU2S3z3UIkxoORMFUe8qwSJHR3civQbDlQ
SiwE9NdIe3Xx8iVeqCPQHX8hFeQ1NwKsSNlQ/jyvvxsXQUHh8NicgSxAjjWzKQHT7unKPChRdU18
BqYBFE2l/H1XO8JUlXkPUcubRYbAySuuqsl0JRKbL6nK7TErDMoY+xf2c3LqRFqfCXXH0ma+kQZV
IniD8OxCh/QNlXArzH59xg1nOdmmKRNtBPok3eehoItg+Vzrjh3VfMiN2t6X/3+qs8lKAm6HSzVQ
3Mwt41c9gz0D5vstHFyXKLDnJnakDlt1ICrdn6HeCs8F8oR2C1AaTg1Z5a1YuAUma9/Cue1AyNNc
m58pzBpGC+zu1SUfnNFuX0CQ+C12yNH7DguUfoRRm6YQHj1HwP0lYqdltAARdWSAoxpBZQR7jXwl
SeQaiSMRiAXJ7KXCJjyDiVihh/fwWUuG55d4U20B15/wPWillJytGePc2xsSDWUFRvZV8EDDLXQr
qDH40kLY8OBYyXLyEPm3OxQVra7/uTCNM/C9JEi+/4ywLH4rL+fMyjjoOMlmGwnonPJpONgbzdoY
nfRnsB2OZMrrzwmfE4/AAffbhO2YX0Pxy83zJ2lC0eLA3moFFEN6lIbjiFKciRKmdm+BwidRW0os
tQtFSnQM7Sz3o89OktLOPl+tul86bX5Hpq6pN5a+s4lrLpoSEQIrZtay6YqNSm4SSryArFU0XTfV
0gBSQkEQoUoHgNrC/GlVAkdUlGxoH6IlMh7YeUpbIICqjt3a4tFjFkPW+7ODbDAg932e8V2aPyu2
zHJ1N2sS412b3CfflnzS2inHLwADD6RZt7vXAcmmNAe7i3QP7fo/VyqFiM3betN3RvnKQIsBk0eq
8qpuIrRFw5gA/ELz8Fk0m5yDpDXzuiqPE4omfOh6xiyJKwdXCu84hJf/BIWtGQbT5X3pyXWhzw77
ix2wajYjtLt7xNJqiW9/IRI6X/1V7z/tiSgFbccnLKD0MBgGHb2CrpN5Q73DQJWLUtWKEyVKRIPN
52luBa3Ou0N96eUVGUlVkSzosQZaeBunT2lffcyyEeR02edchrv8O4ScY0H7I6sbYW9GFhnhgpxk
q1TQWGYI21S9hD4UTWg6q5ryB9IsyfauDfWAOFML4RQ88Mc4jw16VxqIS/NM6xdJ5I/DtAA8FIfS
0jbLhtOKf+rPZqhiCHbpOvKT/1YTAWeNw+zW/iDlAIC/sqIh74v0OqCj7TAwBBvY4J5xmnH5Hj4L
7nuB5d20DaxgDDuyZ7pO8OZIeJWjLdWqGsoKPxnFAcbGoaQhHnU4nRdXzmlaUUOu0qutA1eCcjQW
U4NqDFy9XN+KvwQG1KczM2dtPOt6vmc64WXQ/Ymrkz6s3eS7BEpmwy55oIFdqvJbmIvrzuZmnhri
lqrQMrG0XXRemkJfjoXwSqyTx2Qr3OQkIYw9zIQix3labsSEWUf1DLhklBChEPUsAD/C82EcR8lA
CL7YoRONmQS0jMAJrP6kU986z207+DOe47+h7fMYZSzBqIVRiLtt565ENquXbsd4kkGlycbZZ6pb
RxH50MlDctXGgVcJfrNIQzzQ1OgXmKbhxhdRiYzkLpsKZ0z6EHzDKailGcz0S4Wd2Uc8kZkz44O5
zTL+zhGIxmtfdpqAlaKcQTPPKTTpjuYTLYFJL/VGr0/8q0aQgjxBDboPB8uDwoEB00b+5misp9mU
Mn40zo3tHbluir+3o0IbeDB1+a+2emfiwl8v4/aQ2lUwn2LVzhKco1NZrXVFPx9wCnq9Zh4f7+8P
QauGsLyQR2zOEWSW2KHXH2xs5peWjUQ4z4tuJq5H8PCpHeBUwiUT6wAUoOzQboo4U0MG5RAV7ZWN
yBs3MzgTpiHxbA8LuBahE+A+wlNVBoM1hBvEizVUOZmxKNTXQg0aG8uhuW2jbLAvDVLv9Sd+GSTq
fnXsjIQHQikhyn8GIiN/+WHlPzo/dD5CNkUvsXQn22A0ltmlrSV3gWckfhab+XtBEokA2IbArZkr
a4EkZNUx0d6vtA5AEwMtQ5uXQVnRtaSV8vTClf9EUc5rNJAr808aI6NdxE1A379tqEeBrNSxO6Dr
jlatZQS0Bbd0w+3lUGE8ERzzYk30R1/KS2RA6g8dMyEbaYVCfX3pek3lY7yvVYfSZNpMeDtEWVrZ
peFmMo4UQ7oAxF+UdsYH+n8Z2jT9kTKkeivMR5bhTltGaez4II41WvLFka03me2z5o3CwCYBUPdX
2lQ9Rg5oUV+exc3BemzqTN3XLbNmV89AZfxLYhPuQwD9WKUvBsqQgtjTmhSc79/QqlYCutWClsJX
juujsbbOUxDFD8Ugum+XXMl8MaBlqnaPckklkow0nbu4w78+SsfTa7rR/c9AT/2bnm4+yOK4EkoJ
/bEkIbaJfgmSDW2dby36t8gWcJ+RuOWTz7XLYR6QsFADYDB6l3oK6DaoG8zy12dZ8uUGuXw6+6zx
ExIwWoQExVNrf56R1QStlSF3lJIoeph9BQEfkL7KhwRBzzHpwF9BYDf0WGrIpaAsnUj1yv42Qdbw
oQlpyVg5zTUR88wYUOa6STxSkmeog4SZAiDo+V7QVMNsW84ySZ7NGClY1O9qxZ8XHORGtGp40ILA
OJkcMR8IWnyI60p3bQUlwYoMhXb8Holrt8DbgcrhEcD9sZQ+fLDUkcyzJIYx90Fqb9b+0hEFiiG7
7pJLxuO95jbmLpbrCBykIXoxe6MSUdOFBgwZT+teDqw16Ij0DuvTq6m26kRh2os4bt+hAsVlOSNT
RUQ4An/R4W1P5+UgHWJcoeYHptZKT9YA0H9BttiPqeDCoCs+X1I9x7e2o/Yy017XOBvmYI3iwzVD
aOUKi4nCJDlIT0XVywD6Wy9sxBxOZYxWBE/jttqODArujA1LkU/rPNjDsC+WAPyWhIvcVRXy7COh
LQcu3yHeBwLHAdXHOPcfUDobeDkW+0p3/0zXDy+fTYtvD4tEBkA3k8p4WpgM+2voIFe6OvoxtfXn
5077gZUU3SD80uwv+LLkWiUq7d5QZVDccg0G2Iy7xRSACTAS8jLiAsdZPwLR77Hre0uPg8koETls
yTUAIuqDN7F9alg36q13dfC7G3ADhCl7MuRrUntWLtGA6LEUE8Lb1Z4PMDjVMwl4yrt5L63F5jz5
hP5sdW6qgVpbAW+AP3tZUL13XTe/wHVWOWS7+8P6nqzo4dxbJZXZEidh+S9jdH3DaoZU+gxuiSHu
6QvVvRX9TLqvW0ylMOWLWpPD/hEmYZS3UjCqiF7lM+DfL5/5eihft1jvMQgKNDYCdd4zylaj3YLc
SHG7JJB55qbGnN2agUtKWOxiR1XRBvgPycA5gtqY+zEnOiHzYuUqAw22JdZOzu2QA+RpnZ389qcn
krFJ6EiTg6gV6nPluA6MHvYLz6jWtI/WJuX5G2Us3AkPUJ9WeVoCmkAMLQJXu4EiEJ4M/q0u8q2v
wTdCYcO4WnpB1i6Akhkn6lr9u2peZQZwreWJcgKtiDC0EmfCBU+B4n9wtrWHdkfihg5AiIyepUoD
L6EFbBL6bwFnzrszc5zYX9Qcv9XH22dkparh74Ck/T/XDmbPqU+d1jU8E+FvAZR9wLVk58VZFWTN
HvdyrLSpV8MoxR7F+bPwwFZPn6mHfTqsoq2XxjK1wVAAWJgIPJxvo1xzh/rBUfFniTUxYN6QNQTL
Ds5BNVNLEu7uXoW2Vw/DJ+tcGxxH6Ars9EfJ6BgwgNjyCUjStVXlGINM9M7UBffFnp0amevk+3HQ
w8NSyeBMZSVtZfljJfBYJgd0DUclFGgsr8r7ZMl5zWOBgyIOpbq4qOs6BLO1hzO13TKY0XQA3++H
0yxfNjdpZgrgzUEf1HFvGUmNJo4HprkiFcv5ZXkXrk6sj3dpK30bHKfaJwEuDzoAoUAsGrgkgOhS
tGwIUtdX/92DCgQf2f6RSJebUOvKTKmVon48Fut7ivDeNG3x5uAP/s4eypk5zf6jLULi/cDPyzU3
2c6sk+8QzNMSjM4VAI3N1k0M/WlqulO/SMvT6FFZfr/B2Jp3mlUpBrjMWzm42bE0LC6HcuefXHZP
SfqWhT96RQTCqvEK8HkTMkNiKqa/Fk7DlVzRCfN7a0B+x5rUfjWku4w+rIkfa4CKAecj6KZQ/XR0
ZgPNxoC3fhft03pC+aZuYcejyV/tyaEv1oM6MqgV3Qu8KopVBXyqpTRU7GVjaYQBWaC1Z1V4keEh
YSFyw0Aft+RGyUz7BXAURNBr8/ykSNUMlb0hWWIpqxPnVMN0nNMUE5stUpUsJHKG5OFS3pjxojEB
AIKJwgQXpRm4Hxil3NVf87kIXU4xDBn9e9x+YRBAGILbZVpNI5a3Qqo+hU7jOhRhBWGEIdn4R47V
3pWF5PjjtGAKpq+J3Ww/dpt7t89CM8F7M0zsDoNymSk10xvuOs7eUCzy6telzwBgvSSh14jKvR40
2aY1HiqYkqCTAr7bLlbTj/goMAEsH6EdlvQ/P3cBsQyJnvTnESOEryyaTMZ+hTkA4vA8vE+DQLnu
nsbRHjnd+8lBwtZK/nr/HoWqPPMiFbub6ZlcczouR/KoYWBeHRIcwoJD6Hop+qWzU8eFp+6wRO18
50V58HatKeHpmG/jmrfBJCsDRFLBWaWFOKtqhrnudTlRtWaX65hdOyEp5Oxc9lTavuGnezAyG02H
6swQRE/vz/cmupnr4I6xrj1bqkZnWO4dyuasyhBohtpdunIpcQpBmyVZ2ddljr4lqyBvXR3+fESG
7Cw2glSaOmqqudOhIVgLnt/3GRBFDiwRIgxo3euW98ZzLlCPZjXh8t9MCx4o5G1xEbbIO6+VY092
PEuCLNT/Jo+sVk5XOTaThFP5nLKxtgUOeouupfhbBTABRZOBR6wHHuXQm6T8dGXAl4x9RFchmRS0
QJd2yYhsOQUX+YKAX7orBJ4o8ZSp5dfxqdinxWdPns2NnkWakXVBZY1IFssWO7bqRZapr1hcmoFm
OjUI+Q2fF2bPNlITv4dz++oyzEthsZ9oYh2Uoq94r5OX5hzgyVkQq2nYUrh8hqutAkKWSRtGX8wa
IZOS7DwcwDc4xEgFJvddpnO+XfqCJeYsA8Fv6yzvdrBfm2S8UQz/XGgYIUD3gw1oOmKLNb0+DvWK
JnwY5i/Swho9ZoOeRuh3jDbzxD5zlgznjSjdWzIfUpTyEn/6qOXh0LYy7Di1cLd/eXqFCGNgaCdE
64+udbgnJ3rS3yuN02R0vL9YD+rsgJYYCym8kbUkm9LGzuJwgMi+PLGbKCmbieuYO4MiOi+SgOU7
jWwTbxKNwMtsD1XvH53DTVOM83cl2jHGm9reQdEg0IxG3dfA1/4skWiX3LPTt2GZkqt7qyvTN+yB
q+N+JMJ+1XaJFeI6gZ6WExjozmpDDrc3NujuGIpARhiIKORrm8grb6xXWbRdDSCKYncePjew48qw
xisNsNTJMDtOw8avWNRjF/zxDXqzFIMcFNXzlmt4mIBIeSnBk8XJRzhxS2qF5JVZyHcMLtGF4GRb
4Pfg4KuDG1X1FtZaVRuEfmpmVpqW9Z5ZsA9218cq4j6kpDcOGcnclri/oDBPeoMU+cI6hgY2oaM3
1n+/r65EihpveqpvHd8Zlsbrmtz5ur+tU+30Kx8PnkE44Bcwuev0MseeL2MeVOZyxnKf0UJa0qAy
vlBk+qhUvyZoKcK11+K0g01kYQc7Vc9OVfF8wC5hp1d0uOyGz9BEq3YVJ7tIYt5qH8qrJuuVPDf7
XlEDJRsqgfy2zQJNlWbz6ib93VQsSgLn7rlcnYQ5jlg/bfw6Lv/WOj6eCqfq/h/fgDayU01tXUIf
YJvXJU1W+YNuVYiyI0uPEQUY1ICVQNC2HLg8mqSA2+5JSkp3/dflH50QvpdUWeRt80GNPz6CkhTF
BnRyqiLXV1ohWitP8B5zw4mW0tA7UAwroXQLzmiHMiAvGCOAarltYNJuURSl2hyj6sYN/DWqdZPq
OdfWhkRhiNoR569eG36U0cKj4O4PNAq34GNyhzTR1/+uZ7Krnl/xQQQPrZFQnrN0GLlFUr4UWTYd
A1BNOnf7Exg0lJvpO5fWWH6b7XpkL+5YQQOUIxRgeUPEF+eg/192ea9VPUuaoTad6CYz5VTY9vek
8vyA1ihTKUI15Zyoz6KJNrJUsBeeVfmxRonOgh9xP2sDYj6t1iNkR3iu63XKiLP5tOnU2Ad4pIN6
6gLpuGTRz7aGI7qrlTXXteAeHDZ0sH57l/iPOAy4vg91yFFZSUVIE+4ywmYaE02my4QAtRZ64zFN
S5J+PyYjfwvX9V/O+4P52W6A6Zv9O5NeFKzbDBnGFtUD795i+gFhphazBmnt6ttWrOXU3atHOeG4
dzJS//bdpW55hvC2UFP5DUtMiroq6FMD2K5f3Pr/L0rEflktWRaASlZtZUlg5yFLQAuOSNBgxJHr
4ec9x4b6+xrnETgeTNVzGc95QAFCjOR/yPHhBOyr2XnPZCyAdaeqHgys2IR0hQTmdeSk+WEmFept
PDR4zv5yULpKc0dQSDS7BqO8NRPvpzRNX1JRFLAemdecLtlieHpFmZ9z9z8YzilfDQUUwoJBOnHj
6RnRSM7UAsB1M4xlxQlGsXYcS3os4KHgsgLXdfpNx9ZCksI8t4x/WY+e9PKJnFMmrpAHLTbXJ74I
+5brlAB0H2Ua7W7JTfJh2+flp1GufuFKusjX4uoickVQCuI5rrH6+LuYwjYwJul15m3YXWZQQ9qX
mNvCS6OPQleSfbKaJd4SqVylfptvjuLuSiQc5v0Z3TAqAw1IeO8Xp4IPUZwUM8WyrHUBOZJxo4ML
rfCCEYDlopnoYgSqVcxQcUjtC4vLPXLOMSU78kCnYjiwkfPu+1Td/gpV59NyWcR5ZJ5qAzdSimOO
Rl4G1SpqhTvlgqnd63o9ADgdSVH9qM2OINaSZtUGEuuX+5k4HQuz6ug8CmJBcSZy1gKpTgs+S37e
oBdkwHnNawTm4qdLX/IzooumSJyPzpePXY0ndRx01fr563pYLmkYF0cSc2wKAF4HaDmfh5bJKZyd
eVXFdGYBWmrWwv1Btw31lc910n4qsj+m1+bucTXbhRYVuK+aAPz0Z8VxtOgPd2p8fSbDqAs6tUPx
Y0sO0hbIlMj6BodyzHuwCqwoCjEv183+uFHgurzqeKQGBgjeZveoGhiIz6dOzmAjFoTULx5rVJAZ
/ADcWsSOo5B61WOWkiOvXV9aD4nYnP+xdQv8hwOka8kSlLp7qrbRWCxoAgmUAKNsryey1/nndql+
xcJVl/NJsF9MO1MDh1e4DFtSy24HmFofjTdtGzcqIgDOSlezk0i0iod14tKWaTgJDr63dXZExLW1
Y262anGsyjtXvWnv8xZtH6rVVK5G/BZXF2PcJ+Cm/DAN4of31iiSQng1eT5WKtns4OcquzEzqs2a
okuzV+XobDUUIMOl3KZfKpcgieCaGQhls6gx9oH2i2GzSSN4JtjHkaYBAXHhWcI0Lq0DAlhEJjPj
hLQRplHgatZCNOvLlEnoK82Onx7MSJdxNKa7EKBCRTeYZf/vY00CtgJUaLuSqCN/XLL4JApPRWQG
SgcQFrbJNjQ+XZgTVH8M9AYojFY6g0LC4VeLTbpLvjgxI5CbswBWeu4fs4rFRdw88zNF7PTVDtub
Tla3xffSg9oV5dr7Zo16ijc8jUUK8l3SEZUkVBGprGuhgqqL7noO1/wPm52eowrg5+wKX0+v74Hu
QnoVPVRc2r/KMkRbnu+r7m5LdVyMQhF6OWCPWCSq9ug8zR6kdKAnd40mL7KzHqCJ6BEpzncCycvq
eVtEP/xNN9ZI1p/gALySO3C4wYtrqfsZzhYwmDhpEZtNJZmmmbYEbucIkQYiBErIemkbvl8DV0LI
y20vF2hJ1k9etaIhtg1s0wm5hvlQ+MUq0VnAmqq0XIKyQGKMF0AO0xXYCaDy5rZ+Z2wkv8I4Sy2a
m//4Ct6ZLRUzEJtWL7T8zT+J/C0uVpz0ibXpQv897NpMf/Q0iRVp0rKsY+zzHoYAQ1KmSzumuew4
0n9sPeE+Agidg2SUF6UWPVb31t4jimARzRtjrRFaE/ieACjUQF9x4QBdRjQMzDnbLtkl2zMTkYKR
SX9KAi9rcO3j6Izwlnv4RrhqMHD9PdvivK3arIA2W0YVolW11QzOx9fUYVVu4jcgkAKZzvkc9LTa
+B7ePdlr+/3m9nQ9S1ARidYAVg7Yn6Zhxx+uUwFv93I6wREH3/PcyzFdfGAGLmlRWEY2dXDsln5E
T6DtWURbOg5RoxrqiQ4yFUR8vR1Fke0ESGet39oWTBhm9lrzf1Eznmym1AYLRMJknEQvLX7Vpy06
Z5hBNIu8X7lgDIzkGjUUSM3eFf07dCQndr4c2ol2Ksm2IO6NtK36F5HWQOC6bVJb9b05lxe9llIS
laa13MhJ2Kb8xpbJNX9vfr+mnZ1Wssd3ysLZ+FFPKkAyO+n6mplzhFYqHz/+KbuZueDVxddGzztM
Zh3H4Js9o3dt1f+tybLj4lDlRrmRAYwBwaoMPWkIdKB6KsduD6GL5PXLdkbGEj73StiL5wOzmZNY
ah9e7MVYlZNlTkXBlkrI2/pow86lxWV2JC8n5uFbEDReWtOB5/1LPs9wrJbLnTZscCgVf7gbqOZd
IbqBzQ8j5ZzQKH9EsFpm+CAFo5KAaaJnh3SA3myL8W4FOQ7ov7doaMOLWQ1Zpcy/rjoDdqBlm4UE
qpxfUoIjdg/uSSLNbh/nnsI/ktFv6o5d1nY+VlEri0HSImOslR5eJRoBn+ix5jc2W/mE0yw5WKZU
P7Wo3A/hj+Y8WmouFB5IUw1JfPDjFhzo+XYLoGf6/ydQLVa+WBrNztOWyA/9TQN+6oUjDuOrOG77
PjBIZzTFsErnIEXCwSOOoJaUb8pMDpBvjY6jlaAFVrz6Q4jIvZWP+3FkgA3JI2sTw9dBQQ0DA0JD
igcggff8qVgAtTsKD4xFwWd35gbdOWSWvPQp2geU0rDApaNP07U2LjQMWT97BCV6XbuFYHldbNJH
BBShG7siTjSL8pDVteoSAaYNVkJpX4O+rn6P+qMuAPsZpyBdLEwP0O1nANG6fsDl/DHbKzNb65AA
JVgHTeoZPbd3dQLAYxq7xBQg+4RXb2EEFBrDe/F85vy2eJV/hoWeJe2+EF77l/lTa03milBsxbmT
4WElTla3IFkn5k0T5ArHtGOV4h5B8vwA8TkZNVUN82Rt1oDuxIN+3C5iwKNxraag9aHtQ82VzxIq
nfYX7gji0sd7khezP+IpgPPnPr4XbdPMnHOe1hk7UhlKMHLngMiO/XNGCc0kW5zs2fMYtm6yOuGf
RLN+dJunZdvPOAm70BBJcdUnF3l/sGaTpeFXik3fyOYx4VdeoiHQEmor5rDKWVD1YyhCEUv4AkjI
nyRI6s4O9I9FCzigPCsAgpcT5TXCMyj9rT4h7FCi6w4iuUkqAOThtdv66xtoLhEmQIVvbMcSbBKK
eESQiOpjTBWLo6IiqCbquEAqTquXA/VVWUcdwWDy8QmlLuvuBXub8uikgawfSKla7/faIBqDsw+4
SPzMMlb8aSZGtShRC+uIf1SvgVsCTnKgTbxwFZ9LmH9HbDJuC2ccBgt1JIg6/ukMOheuFfwaT2l6
03WV+BRx+PnPnbx4eMwn2OvDkGTZAp9tO3G8QcUMbm2/OVAd97MtKY7uwMCJeBeB14LoM7OUxB3u
T7W3iep4tgomTq29xUrHtpmxM8alF+kWEv18RWHLPEmDR6YMKu5Ell2dTpBaiJhkOZScoe7jn472
C+jIBawHGi18hDhnvT55sHvYKSVwJlCaTiLjSAu91OM+rNOhE9GRAUuQyjpWewuVZyyoHzYXbzQy
3cRYn4Hb3VbdyQd3Zj+NI9aKWPGvubnOPvIXmSNSgcDpjDfafphXeyRMZcdd/7+f9rEucTRqo+d3
C/hZbCZkLqDYH3VbOctjuorPAC3537OTM9huBFyEzMcj9oo7kJxWWzRk6PB2HLHnnhJpZd1yrgRT
HDLRo/WXN5GAVbkudqz+k2j1c0Mbu91RoV6wcauWZxTyUp7eBrwc5B3/5iqcoXasrpbvlJA5GX5Q
xbvxB509+Q6z0BboXjDFJKymVpMazeFOc+OC09FeGbwbvMtBTXm8IvnzooPPEugqI/zcpYwoojje
biqmrCqNJutRg+xHo6fD976uMYxY/9Ikhyv9djkJskXPuLmGSeEqExqnBs1eQygS2c7lD4+UiWWr
UtJJlu5BGk4kMxIVf7Dn04iWKuSLcnwU1fhwBb273hkwDUk8UatdfcbUdXMcgtdMEMAj8pRieKa3
l0oTahhSyRxuZlEvbwj1/UICUa+zItbb+DcLsfPEorGI5midJb6AX81/RdxXEUeZFSjCLniaajzu
uGedRekPqWxY8e74D0MVgKIxn56cUSuk6YUTDznYWe1aqnvPlRyviVDbYj65sNkySchl1+kHUIeU
YsNPBUrqzWBjKOE4+OuU/eTtXoRxrMwFetzNuWQdw7e01Qru5cRfpZzrTyT8GxcDDNUmCV/tf4v/
45iIuwj84V6uLR/5QTpdiSG4CmgNq0HZW74rDTGeDzVtvOdxMnS4DMW4zHlLuhQMgs/f39PVd/BC
kL20pLbcxbw7XXlIWWx9Ij0PqfVkcbSlbZplq7GMXfA6oKyooakZBjz0MvkcH4yD938/IzBP0kXL
e6H5xOvc9gggLA/5ArxVHrhHcAatqN45szzwUxDJ55Jp+djVLXHcHVyLrT8xyUGtntZDZACvpSf1
UpAPLufLsnq2hJc2+FvxoV2NUyEsk/MoG/V033RpX7vZCmQb7Mix/LJtwt/AuKtHpPubxOJY57OM
xNUzNWd52ifOGh0v16RlxxvI0c1w8D2907rF26gBxM+z/cbJ55sP5HY0XvYxhS8dkkSQs5zpRB/e
MX00RzAa++eUZkKxhxm4xN7a8P8oBWa9EswekeCcixcjxYKPBr4UpzPDYxoDryYXftNDtmbitV8I
bL6E3WQHhO/O92AcmPHcqlOj5zkRGWvl0oNCZ2Kc1W/uE3GsUgrNTWWLtbJNt/bMO87KSSAdrwrF
+9b77rABq4Zoxtb9HYTLbcM1xFk//V+kpa1CcK83ecdMWWkYh7/WdtWyvCI9YHIhKs34cuGuKkFv
rlS2RbBFdWabwHybnGKlLxPiROlBv5ai10PuRWY9TlEaPgBaurpE+/7Zr5yzlmtXwm9j9j0eSt8v
Dg3IUuoe/bRPOrtq2yXlJqIkIMZh8TULZbPWFiGPc4Xm4++dPXzv9uU8wkyVsfX00nfXPFW2+m+E
hEexwIeYDtpHJ7oMstwjhPzht8n+S7UJ0qGJZjks6LMXoXYlbZFmwdDoCJjzW8sKaWR/ZaXnerlW
knroGFUZEorRGTOpYI9rEL1zMR/zgOxqhc1lOxXyM0mMgqBHZtycdhpJ9JUk98mg+WTZ2PWl9bxx
B6/UcvaU8gGTNZUWy2roVBCfOrss0pTc5eu3jpqYekey6xyP55wVCg13rUbg2vMMLvtt2biJI88j
ATb4a7OZT9p2pcET+uNCEO/MnM4rWRqsswSVUCWPgy/gR7Q7qdEUiwPTGcS0bgWQobl1d7TgAvyu
2PSr4DCdNmEQTIb6crFPlyIVOjPzM9szVkIIeGCysd9L/nWxb1w6VIGi7CCNDozVVEZviWL8LhBv
mlc0H7ubhmQKM3KJyiku5PyEn1Zal78a4MUetoXfQ5BNG+dZ5A6JYsGbvvtgNoKZ0z+A1U4GA4bF
+J4+49U7VzTd69ZnWhvkWL1Y29E2vQtP/ogcZSgWDHPCBA8DBl+h6IIDEX3df6iTcBrSYfWynCYH
d9bihXEuuksffay/2fUdZVD2JH7J+f3BqTkuAGEU+PmeuTY+ijKa0W1G8OJB1XIMmelkQsd6dCQH
a4uwYoD845KbBP4cMV26sxyVQYPO4cYYNGDix+NA1raTJEP3O29MF4Q4FtRyKRyE0v/Bl9X5wctQ
Rni7QeiFDWiaJKoAscS+dlqcd66pvbH4O5v/HfwS5+sKmVh+1ZLrrHV8bkq/v53t7J1LFlxdzWVh
xtr4LALsP0xOEx82jF3AYg2QhPFYhdjPdfBdOvOhcbDLzitQZBZMLglvonKEfTkf5glbgqeowLSQ
L8YvFn/ksuxmxqS0ClSsj56ar63Sri+rBnfXdWxWSDzECyr8ziNuUllRLt/sYi9NYfs5ODjYHtcn
02srJEWjXEBZ8l6hddwA3C/UaoHTsgnIieSjJ7YYpN1y+dtGkgbHTwMxxFO2i94h7XfzZVUuZqjE
GwZSqbQF/3lNAmUGQ8mV7SG9nKgc0pXWAjXZWLEvXmSjG464QoCKG+Cdd9OBtsuXYSAIzlyujxq6
u+SvZxyBGfTqqUvN3kh1wcmNlZHJZ++/OaeNzRgCKAuI2SttEUjFMm37HZ1vTaxQiBk11SsWKHZA
xJogMt2giO3aWspFK1tuqfpujMTjYVZU8TdHEtR6YAdsUxhd/IcS9/QkaHaCVPO1CXC5HrGg3JNp
DmkkBU2ObJ++5YWyNrlALAukOBmTTJmJbYdiD11LhMr3jxGfunpaQJjcpikht8ZpJ0VzIfRgcSyo
7wLqmCKKOTeD+ZK3d8+/b1mBm2AeZAL7GY7K0CWadaxR7cbXEOA5nbZV+8u7rQMmgCl4QKh9Bkeq
NO+09ss33fQ4Dq+2aeiAgeCLjpTD/oI/Ft+8V1xpvVhLDQsAv7ovlud1HVfpiFnFn24LxJv1Mr8n
A8/awxRAJEuYSGAPvcFkNJ2yzfcHp8UiAl8yem9eoVLScs/B8LcE6HnhsWxeDdzIgoqqKCPjaSdf
D2D4OvSaFQHmEdsNrFq+IYXIGKKI4B6fL7q5booQ9ndj/uHjGwEWwBqErqxPuJe00pTIqx8A6iG2
i/u2E5iy8GXvQhG32qV4qPTsfZTl+YwEd42RlyGjakhQsL3DTeEoYEAd1v/ROtfg1zX4nUaPadnU
JPTrQQi+x/1xCz6wyu1RjdbI04yXXtXiShPOWfNjMUqEKQK9qHmV57sXe42vviRsph2/Nb5zTN1W
qoufg6RYi1MVp4iiju84dvV/9djv4MeK8ZB381Cl+GC/WIQL9dFtkLouKv7N2kILmVKDsYReH8hr
n6hQHqEaASN4rcpl0v1ETowDYq5wi/VCIK38YddS09hPgW5fjDJFcDU4OjjOIlAbwCQrj1tm8GSv
RBNkRDPj9zcedZwKFkBQp5gPHdv/bOfRfx2JQ10Q1CRH7bjzrKR7G4sl8mg/NVHUQ/25g+dfIFNz
fWvpX6vZwr2I4F4tC1z9ZP8DI+456xFTP66IYPQAHVF6O2IdB6kEVl/l/heJlou0qednvTgUsCCW
XFhSQeFi54wbfyettrmAJbtsHAh6H9G4JLpKn+5IbAHl4BPgC9SQv4GUxsGSt+Y24WVdSrI/IDRl
flE5gUm8BO748N8R+7kCnGnNFjOJ0yMpB35nd3KPQ35PX145tN5j7grS8J2FPBZTHavHvoVzT/4J
zAcPviChD7IXDoHd64MMIbJmxkVTsPm6fWstTJp00lKHdfnKOe3mQG/yn87fKQnIJ/WooqpI9LlS
rnpTZcxEyGyvlrmgU4E4ijyjBAKjTl7csSdVFdqFiGOhmx9vEammF1/PXJNIwpp/KrBKxwBHPhdh
o1BsqP8mAKYlsjEZQsLs58q9c5jNtAhlygPuJ6lRLMI0BWzDtdxNuNCUd4D4GGiTndEoy+dxW2cH
L16FkvCq9M+4aGFAHPfXawQ0rJyzcqFLAB41po69TAovExJR4lSi/NZXMLz1RTiGOfWI0Ipf1fzr
tYZcC8jbPIm1TAaTTjJcz6wpmCYUq9g/c0V3hq9AU747a8T7uggWTWAUC6XfSp+68OcLsxBfKUKG
9lGxx9Y3bsMCAuPJy5lX3MXj8h8H4tyCLhBCU9PzE19a8mWzhZJYQJCTKBfR26GIpAEZ4E0SPCtk
vHnr9wuWfu9mnB8ejz0Thmksvb2kUP/SRClaMu8mAqtoCZzcFNq3wkF9G6vTiEyNIoC7UzyJLgnx
UmPJ/Xn6ShnVx/1rFw1avV4OMCnvdVb3qNYfSCvHChXgZuZbcHa01D+JuT8QxOXSTHP8/hk5QYjy
Tp5KkSLN5kqOcl8PxJxwz+1L/u1qfCwT1+PU2FcLq+gUz33zJ7OGx35pUyZzLBvr3s6SMtUZSwUo
Th/ZVezjNQEfHKWz5W8ba+v96TC5kB+94HxgmohdpppCS7yTQm6GR1uhu33mP3CdOooP9lwqB4+d
bB/5gahsl/wSB6Sy+Fqkncb5wqqy/JOEu0rWetBmxjJ0tLluAIJmrESy6xyJzc9xHh8JOJt+oHyH
oQHC4ucjJTV6LRTyXfPpg2Nmzm6T0cWI6AQfdKOut1iDYoi1hpjBX4nnc8kgOALo4BfTT0EQFqY/
/mx5+Eavq93aqmUWSvwgoaOU5G/umqVljhnRJjqOy4X667lFWfLh+jGgMBl331AC2rz5Tb9jp3E0
ZWhi07bkHr+o2dJ+nl6NEdQHtzaSu9xisHGiSIIh2mfIvLVLlCxLqH2Z868sn+iYsl1YHTCd08wF
Scm9MKY4MA4gZTgWyq97prvTXpxNj+YXKFDtvcAGblyilE2hDGuj/I7DzI94wCq/uIP0vz8utOXu
EN9Vix+DuWYaAKsLXFn6bdkq13gQuFjEGcLjQOi4L0tQALBC/N3QKvIpH1zKFZi/5scrVtxWrq2g
jDwBv3j4GU/4KVJaYVOwN7/In3eQiZj2UKxT1s/8UMSLpxN3+rOUGvoes4ULNK91rhwDOU07c31G
GYkM1Zj7RczC/qOgExiP6vBvcz6ihD1QrI4b9edLZXBWPLdn8HJWlOUTl1bMsmxLeW5KaCdUQrvL
R3l8TnQ9IFFFcMaXzmmUvYpdFMFsf5joXns5oAVJ5vfddyAQVIpSav8nxBgvEXBv5CALXC4ltIyB
kb9gF4B5U+VYn8PbO1P7Sl47FVnXxaHgc9YYpBaPa/JIbjgxcdyMBdw78kFCbEJYpIBIYMoZtvUy
V/tU3OCQMhNSWvEWvNdo6dJsqhYLcM0OlX0ktBATEDo84Detuhxazu5/uvj6xPcjwEOYSHffD41a
+bjSVrwTQk9FHhSlEgd6z4Wlh3v8T3PvHw76nbEQ0S9YMY16yw5iuGUwYtpehtALOSrrFAKgr/nQ
3Z7oEb5ii3sW20ySqv7S4Z5nfA6EFypIBen/3dOonJZRQOp9nhVrfdY/2caQTZ3lRNnTe6GThO+2
sBGwk55eNDE6C5vtF7sWS1Nc7NqjikFs8LkUqfBAD+iIiCsKLZoIg8VswjW9Ru8zbxtgJBS9Oowa
8h4jxw4WA8dtnrfdse/DMzX22+SieBINh3w8KeY1+cvyrHL3MRoHpUOWKYgEddF/EfHvtN1sZqMZ
aG2hD9M6JMOV4nfmttFbVxJw4/9TYBJmvsC2E6eLX8ny9TgjHv0c8/pTLJsFI2t73ut8FmNqNOqY
91o9IPwppczUQEMNLkrjH1H8MDe1Srx+yayj7khfvW3pqSx1ASYleVJA4TJJgc0afXoWk9uaYN18
NprvNRMqEGqhZR45Js+kdnGwtvm/rPrz9Dx+jIKmsRPilpzkvVdd2MgZ508qQW8wt95yQnnhMcW9
NP+7qYgJM6Ny4mV1UewqB1LOEWRNhqM+suRtg9bFSJVEh+86rmBCO69u6HpYxTuhWKqv4yaHUeRd
ODeEiTezoIotiPcKWs/ADbl6zgdiG/SYWQPMFWGtYI/5y1D0LPS6st7onOyqtiDsAD4/bgqOgvXu
OAsbJvce0Jr3+DkN61ON96k3ybIzpjQ5bCdEOiyxEbP8J9BB166BFb5aURReKBtpWR29/5R0A4iI
1GWK2tJw4+l3s01CKTqGs1B84hNXM3ztQlLGwKjBK3uGRwd0ajLyqjix4hiFfOqgQAvamHR4PF3P
R5lj6D9PKLRom139w6AM5pZiymlG6r5QSnkHdBTV4weL6ufH2flB/GzrIb47XZ2k9j2t1WP5Kg5z
MoJhn2dz5N1n2e4F6iOJkbCyqZVDqwXsYqOMoXhh3ugjr8a5V4zcmWVg32zjn2wH9USecU8eubZ4
NzpcRAC74zzWQueCE10WG70x8rmW+oNs0bZFzRffIc5yck/GkX/Qzjn6dcOcQ1cBEG3KE2ZymMJd
+oIjv+CRA4dhnlbOytoB4aaPM/cFdSgkWzir5zTEq8VVn7/9nGNJOusr1c3OGvqftpc7x7PZLEOD
DE3isETCyEuBWm/wR0WSKgR2cGbLiKva58ELHcV8iRGAQpw5Bh8pxLco9KT4xN+8ZMiSXhF+v15M
n2occ9/TTmMF1+JAsU5FvgNNRoUMStRyl7Kd2l9gju9nGxrSaH8EB8Bhx61J6Ag/1H8xmDZBTuFa
brkoRXmBDz7AOiDjlTB21nyTcdvIHnKvYs5cYAqRagB72iOz4l9w4UGP1i6eky4lZB7oljhaIPY/
+cTDNuxMp2dwcpSE3lL2EydZ0xtspIcOR3GbK6Eomz1+qRI/GB1+6LzwgfqzMWvVdfBIyfNg4bqW
ULnXylQt6KA3ILqsaBGj90Ux3zm4N3o4OtA4XMQmNK6IO6b/CzJR2WMsqeh5NmLW0ha4b+OX+b/x
FRzYO68GBVa+Q3rDl974LnUVBzKu5lJgQcC5gYqnVutHGKlzoByvzbwuoiNC6cxuZ1RSuydPAFFH
R5Ep8YiVsQUgnlyUgHrJata/haKu7G+wAlwR4+bWrN7+frBRs8yFJ9jfmnuCzJCFpPhoIS3TBM8X
xT0OZaKvE/MAJDnDn58dQcxDQNMA02RyHZfbmVmYbqvLj+f/5of254j6sRCdYItyUFu6NZKAogb4
3W4aFC5SAC078i3RqOMwM7kilHuEqYa10PwhZ2c8qy/iQSlzZfAp/c5mdkIlFe4k4P6iBGgBJfPv
LZyy17zLaGDJIh/QLSW6jncW883IUcCUvPfoT8/AWYNg99hS0het6Voqrvf/dO8yPOMedQbbqRrX
G0/J21rcI5+EDL8gac7wy2hLJ0eD6bNXvJvqDmpbfCMYbdXpdt6h/viWek1N20uIDDZwkqz4vBmP
i7XygQgp1ClJAcCEptsGsVYa9dmJGXt/bCCqkHUAUk8/FPBD2JOpQ+akpp8aKrT8cH0u88WxAWdV
bGEbFEe+13/3TA3LbUy4KDA+N0UU3cYyKepg7AE0bO7DmyIfcFGdUZkl+vt59rtPCl+1Yec3SZP8
jZo7XSxA3QX762codWhAsmUAVof1dTzbECrySzPAMh+cjVFAe/VAeOpVlMv5P0ZE36Wt5qbYw7sP
GVtYfC65Xo35uT07pabUzSZvLdfzL0oBmZNnoLrOmYVyUah/52P5xoS8ZgcloFKXf1k23/JZNgx5
AC0c5PP0266tzk3+zq7u9uqyP9i+uaeUt52jh5Xw4r4WGJftYePKOqvS2VPRakXlsWt6Rtw8GSFq
HULK/XXrhnJMtX2v6+0hdZb28XN5kGOvpAbf9eC0z0kpBk0zD5EtAPKxppCWkqFo/Jh7E9zQH9lp
Zgynyib6oWwqrtOFI+aGFObz21bXBJVmae8BWomr84ytTu7ltYIC6X+fs50H2++zipy8lloZU9J9
O9GADyueeauT6evdSCWxD22GGvcyQVb7D7F6LE7EPMJQVik0euuek4mSMjkkjPJSC1iL4ztP/pMp
AS4ctPqmIpxr2s0XogR4M49Arm64498wKzm0xcLO8m7OGb5rWna8hOukVdrP4OFgocvUJ9kSGdYP
H9lFALRcfb3jfKXOF/QD2EdSBnEtW8m9QY3qxFZrETle0qg9xaUlaeAHqHB8afDracdWpIymbLTX
omUeqLJlffSYhSE8mb11pRUS5CXgXWfAdQyJNDdKQwR+M5MmcjKCd2dsYYw9wIu11aeJCEWoDBYl
HE2MATN51C2zfCcLnxNIqQd5gYmbgJDDDKXx+ucZYsE8SBXnhkKCz7N3XgIKaKxFX9LIdW9ZPPGH
/Vm+4jJPhhTTeIhXNvQRH7w4QhG1np+kV34U0kjhUx7ujdtpM8s8s7FyG9O+hdjmoRZ2nRissX+3
PFMmU4fJSXahq/IRh4pcuvr7dS9LVPLj0uJLATidpPOqaRIf/k7Upzqnzvh3/bPxjrLUoAkkXPF8
FbUV+n6Yru9YleAgMEB2STdz5yJLxD/2fWCN9K4iUlmjZBESgGUuRjKZlZ6Do8OJQ1DqCgoU/Ohx
RHNzulzeBlP43O3sGjXcVHYDlPiuqvCyIWRGunGK4dkAs6Wg0P1NIXWzR1T+5xCbMB6vWk92Nwv2
/cF3+LL9clNa6U+E+G6o18Vh/hg27PTqV9UgqZmB1rW4Krw135JxHkfy4MW3TOwim3W1ia7i6KiX
m+UcSMEDFROYDJitLXdgmUgzVAAHhSWuocA+s5Bz+yzbeTWZkKQz3JYFJ6fb4GuJRNaCdtKzLCkV
i7msPyOvitAG9gmqA02u3ykJKc8fyLmOehQOTahmSzzhGUNJEaZY8uPqKYz5rRGi36gdroIIrrtA
ginbCp5+h83v3gmCeLJp+J5E+zt7UFj9S3YnV4A2XF9gfPM+hWDR1ss1g9B26l3PZtH3EnF4Nl1c
pDQERhSQuIknJUDcWeIrA78BQVa9NnaxC0VRN243B2lvoafoiVgr28i9jrVHjjvgFVnjzkGHQb44
0XigwrugY3X+16Rm63qhfo6OdBCHRQqA13+ITLXa67uTISwHq+ywQM1YNN1yyqaI8KA8u3SONuD1
T5EU0eETVHrOd8z8Sz5+YYR/vexNEkkBzEuFE+j1giHRXr3chL0dj64NiJRD1ke3GbWro9rwGnbn
mViPh7xfcIhHHp6Tss9q8us+rjnIrJKfMExdETdgfTcL60lR6wNr380zmx544A5BZWZRHwA/vnp3
VN4hEZWh42l1P2dhJVYSCDM8m1idoYV1cPCdLCH7r2DhSPl0ww9wxLmVF+ObNGhyC0JbdfnE7HDU
kfPYM4qwk8JrVbb46nAbpljdz88o0HtmuDkzILF2LtpXut82fKF4HKVAUM08ccvQKuLWkTZWEPat
t05b+SHcXX5S77LAUqOCi9XGeJAmZoPcJFnPgHSgweM7/s/MH/DoXUqWewjjrAkhdOMotm9myorr
jxMsccgwLX+nTM2WeSpjzcVMgabbOo6vVGdJAs22ZZFf4Mz+/GB9kNGr9MYBqpqsKf4acw46U+wQ
mr5iYBkX2UQ7XttXErslg84GK9AfP7jBuUZbRe75cHexBUzFdKESW5p5StoLSkXtMBAvKIKHg6E7
NK4Zue92I7tAh9+EFqDpnvWCZS1RFU3zjCB1YIPHGED9VzBeLR33K8BubSiIlJncIeyuOooybR9+
0EpH162VZaZCR1DVYxXCFXzGgT93DMgcKsAVuxUsfM7Jjtw+z+PJcibjIcTgixE+YHl4vrvWiFCt
5VHYm7d/w6K4Nmu0aNOFyTXJuQ4EkM3clHe9QmUPr8fAR/fl+ON3UUuJFCb/OT+bbpioM9KGFSjh
wYfj3ct+2/9PDe6PXmiLZni4SvI/8Rylj7l0GAXJmlfUneWIFX+yrIQce+mXTtTpUEefri7xePtN
dfeqvW3mr2jU69IXPsTOs6c63xWZ2oYiM3XPAJtrV3XCpULD6eejiQUJJhw1aqQk3/41/vs0NC5+
U2w7ONEwcw3iaXf0gdVvOM2GQFJ0LUKzZSrzR3l/Duq27dijLTvHVBTQCWLAm1hMel02STuifsc2
yhZTJ2H1RZsMfFMaZKn2NspgBH1sNezbRdwMJOxMiWngcKPlZOiVReN78TQhm210efMxQ0zi0jBb
H5qnn+KVvY9WDpwvCUsvkA1H+OW87/Iw2zhb8sfLCIcFqV23JXYbi65kCVsh7Dgyd4B6/cv8fGxi
Y69MUZqq6fPv1LfGGmC5zVXEvkxlbCZSmDmJydp/lVHtRKcGDNgT+YRda2l1FP93zHRiujt7xSTH
LVU+Wxe9LZZ3CeukYwE0b9gMO1x2vEyItnBB5n9sWgtx543gvQdtdQqN5XiY6XmwJUvkNDLpCuxN
RITVQDNa8QKrUWke/JTsQGFArvOiSmQM3JK3rqUcEUJ7sWSZJeA1r7NAxyow27XS5r9p40uhNXDo
EySPgiZc382/RG75wq9oBz4s5UvzeV15ce+7aBMP0xWGxR8XfjwAghNMNds5CyhAIwUsRyKu6U2i
m2DZTWAvVgXqADHOdw4LlyziRhPqYsu+fqKbzkyc7N5EUa/ELFozZEfYCu9OfiR+DzJR1LG3m+bq
EHIkD7xmGYk3147L9RqZFTBgd6iyUpcQiplUdz+n7nY8/F8MtBJGVeECBT7raX4RjPmDuNsox0xO
1OnS7n7EFvSslk7C5LucZJCUvP081Bbxud5b5EczRTRdHi6tAiWqDAbUxUSYWg/eSnBKLgJB6555
2SS9099bK2hFx0n+375NK3u76JkD7MdqxHvje3437CVCcfZnTwh4Lh/BYvQmEo4gYuJGPjRPWU8u
0COCIl+dHyu+xFxlZj4SqQSh1DMUD40GS+pV23yMbDn0EggNOfSiCWGAIGaJEDkR7qFGzenyhoYQ
FJnq8CVPrOh4DYx90acGUI33SHkErTXAGKOgKQ5AJU7UCqd1FN/fRTqyuTI5fjmJRfY5L0a7b94X
yvYsU+cxEXG+Q27s5xgaxH3dgEUppvnJBVarYhpiadUbNUf0NhvkR8+Sw327t2/YjPgECOyFYBlS
iXa6KzC4gfjdZPy0lTD4qZu9x/GLQ3X6WrNR1L3f0c7rTOLkd2wE4v16309c+aaFOnMKPJIkofMD
UALu7BQobLKegyx53n81mTFhrjwuwp1vzjMdDJcbUyXx7ia3FvyWlh3E6kKnGlH3wOaZTqZX2Q3z
QxCXvYMbY6DquUWJHhkfUsdl0mjhqw2zcHe90sGdQpN3icg0+HL7n/5EVfI4PeLShN4tOMvAHfC5
tFHqvLKjHll9DjCxQt1gkNyVz28pPzEpFd7r7eizzkZMJFSLnQR/fnF7rorsjFqG4bv3Vuh44a1i
njcJSQUONueejqzfsSbTbS+fD+cXs76i3JEfDe/+MR7c15DmPfN9lxOM605Ne0HZCCK4nkwQ6iyY
o6sgh7WZy6fuA1aGtMyB28Mmdct1SkmARWH8E7ipJ6+5gxAH3Lxccb0iH2ucnACwCc2GDUHGKIZ5
/LE70lIKd1qLRZ0llMUS/zPZ01aQhuAgyZSQtP2CLqPLuNgB1g4+X4s392xqZOxaYAkLAGTKW9hF
qCrNnvNwY/xes2YD+yubsfWyNllVjttOwwuh2MwXkfNfRikLCv3T3tIUFDKx/wiD0584RXhMSqj6
5FDxsCfd0mICdU+1RJJSi5VWXmdsKki3x7ydlEuNBmIa+g7Csjixv7Ks5+HOzpKqQvgnoFWtWsvI
1ehuoEgCaFqtGr5PGPzsdklqqWbyY2RwGZOqUPG6OPPMp7buhKaVwPZIcBjTKDfhp8LmHBLk80Oy
b34Kpt3L1C5GE153riwm7dmIPO1uo6XXZPSaWAClJE1mRfjqxHTo5w9BOT8dKfyZ761jxYH67YHV
euzNK7Ap+yzGaUSKRtqxH4I5Kkf/bxmm3cr17eiq4cFlG4vC4aN1Ii82NaYW/SpY4yuEw9jlumfo
DyZzhnDeefXdBGNUHNRvUW+wJXa+adSXsJ43HpsQUN7LPxijSJdtH842huH+mPZkNrnoSdAQbvtl
FGYL6/JZFViV/rcrkO8mKz3pDULeShMpHMlKqqdn5YE8/i3YExAdGAQPx6hQDZrwcDa3FN4TJHPD
5rhxeQWenrw5bb3BGAckqguVc/mS5u7X2/8n49t1LNLsnWg2rkY6qKF/O/N+JkvDu1cQ5mt9nlvN
b5c1CkToMVenz4fb7c9d0yTgs8Sc8oEsdydYwhHJUCBoC3nHgSeLamZLcZph8u4F7qw7QI+V8d/p
XcAexRmwNqjCg3sxZ6P9eAlO3uC6Q8JT1FtxmEvL9YGGF4fwKiyIe/jZGxFdYBDqT8hGrlo+Bbfv
AppNg1pf1Kg4HIo2tEwwC1Tt1a660uQrOIPZF7FMLjIBs1MrsUYpzc1j8no2Ic+KbhjHAelKveSn
D9EA26v2D/BIDovhFJspP8l0o7WIXpEiEl0PjHEdO+3pWkKtLu97psZAb3JOKlQ1cc5Jr0Vp+J4N
pNRCqt1O8nk8et+srD3vMnZg/X/tj2QWyRQqKvx5Z4JFNYNVikXYyM+8StTtEbzuK1jUWD6xwL9k
HquoqaAseHHOayh/mYBQCjV7awFS2i3KJKELeWT75XrOnV9DhRaQ3XjM/e+alaAWuR1DlF2l90S2
vx8vQfdbR7vm+biiUegOZnQgQJyL+vzLIyi3z6ZNdkTLKQlQUigqJgrN2aflekcUkD9o9fNTMYsY
otr3rwGDo1csZxSwC1Y2Sb6hyVEhDbLr80rt3vKEjgq/pehfX5d2RKEvucYuJFO8a+nNU3z6f57Z
uwY+Ev5ypFADJdHeEwCrYDKsZD5lgbAaGUqL/IGNEdqcDSKkLfqW1f6nWrxq8NAqKv8ZJN8vbEPV
Jx7JSOCf5G2aQtkm5jI2BAUKA8Nwi8rb1MT2DgQtNoZOrQkFRV9XLK5b0Lak0en2MyaJI+gT0tfp
7RmZU78DWBVOJt/xSm/MgenHnSU5Uq9N4SkzXt8/O3OgpGJyklV+Fis3pyh4V/TpIdJGwUMXpunL
jeHrNcBPQZPPENFLIx56B2e4JcOoPA2r9Xasm+lAApFEDrBvpdYnHVN/9TWecEeYD9GWqAJKIOde
xf1t2NUzArZiYoaRA0jIgGDoQZ2OMdcK6C9GdEVkAdbg0DsuQ+N6NLVlPZONaqlSrqkcU8m4Hx/X
iQX6IOkAco8NZQk9gfIaBVrR0K8WxYuBES8JbwMolDI23HmcWTt01s0cEeJ6ktXMxJgdbC2Q0Emi
a2n9aAt9DLoxCCHI9nCqUssKMX2A0Wg7L262nwAAYgN6tP5wDwT+SiAM/o5JpI08TIj72OcDE/Nk
70ow8jz5mptKMDceK2zca8pWDKi3rKR/VdRHVRhgsHn+EGk0w39U/CBQmOQiUrBlyAqUrPHJdiiJ
Svw4uJJqFes7B0oU+jGTx3hPGE+lh+wZCuuFvKvfXiz5dbSU0Qv5fDtehSklTLEg8DXHf9K1HPm4
ndVFr554lBDKZP4kbOlRsEYDnyhfUBzgIMZSW+zbuHbgrjTJMMkEqp5/iCJa8fDU4h4SuwAUAnhv
l4mSt+UBlTjMAPVcSfkC8ocpL43OCUt0d/0Htx9XeQFAtWAM09MP26bR+JA4PDOS2ptf+3JdjZsY
PmqmDz/SjkncKsacX36WC0J3WFgGqzfYcPTg5ORQfoVYAMTxfS/jdVGhwBQBg08/JvyDX3U6rU32
v1aCLXNQydbuNyHDV4yxFVr/Vaftx9Poky2O86qxQhaPYXjkVWjJ51TB5S46Y+LK8ti5ivmSqw30
1dgHQkORcsqibIH75FT47o+bQEHEuno27qA6JSsmVgWS5z0c4tNXasfcUWd+kY0Q4T+PcxkvJYpM
KHZUVXlHb6/0tOtypdEAgLBAmmSpXjpw8jUnxefl/fqua/TZQfkwS8bA/7J4KwiCcRKR5NH9Ysw2
FWQwNmVHP6T+12RaGTUodLKcpLkq2hGEyMqZHLNPoMQkGPntRuRWXIiI0PQHhK41T+gdxYRGjDp5
k5CVFpNP4iJujWJJYFA4AuPo4W8CPt5B6O3opwUA41kBJF43DGc7IisNyZ+G5ruX4EwvDuc+sjH7
ASroqWpv7WFdWIaiu7gKq0xzx0ouFrMzlRqwF+Z5fUCftic4Ho1c5EoqtFlG5PPtUPLE0dS3be5l
Chz65K1YtrV63xDNoQA0rMX5GDguH6KLVrRVVoQOZaX8h7/mV/sv8i01Kuo7Nh2uDM3dM3ehoP+g
RjZ6WI2fgl64WfEflTp37hh2WQsKrtlRYkj2LMtx4EVyYukqlAjlUiwqQwHyQE81sKs4YfnXcM2h
ZgmhkBva4mfSJYbUq13hCT6wvlVApxT0He+2cjGANpeYI6ohqscejwKMweRyPHgaUMblQ/gldbAY
GLm3bNtenhO++3zKBB8gvozsjq/z3xG//uOl+jjslbk4YKG4JRKNRfrfL1zlsU/ZxY7BBOQafyyr
J9eG9fDHey0TPTDFxnqDZyUcsX9PAljRbqcVz86eMU5fS3zqER+My1DjcRgFmqX+NfJf928s+Sj0
dCIDAWnVGObiZN514Z2+eG6QYEIlX6RTJiPybnHrFHAVGQ3adqHMjbzwxPbm1itikKUrYdJdf4DE
/HG05pjRvMKiBiS78HYTX9a8mW71mVIp2wU43tDucyUU2n6nkHsCevqkv3Q1ErgU1FAAnvmGcbPt
uxVEIDskFtfFVSza2ync0nSdlAt7biwW8KG5aXLEqLrRhVk91Q7lemm4p2tEbEbJlOdbEveELYQY
razK96Pmd9qb1Fk8ngvSvT2lx0aANnZWxz/uk6yjQmjxGpo+vzZQSxLVEnEUwsEEqd0r5Zp40uRL
3ydLBd+TknZ4c0FIV+lCkpvpeqLb4w+wmVk2TFxAX5KT6DyILnZDXTrrH7Pg4IpNEoIO0Ta7FcWq
ZxhLUd8dG3V6kabanmyLy1EK2oJ1WSFHFYcXQCYCl4r1K3Ze8dt7NltPmdQqndVkQAkqfaPGdDSr
ei3PPgrcy5laztFKG1C1BA9kYll4paZ2IEIm7l2aiwVThVFWQbW6W4PGk8yMLhO7Oa618WlvQmy3
NPVrjOKL2Tu1OCuWNHmrGaQiFp5GbS8VgW4sJUf5tJCUXqM+fSXfx7GI/r16pAgRhn3rCr94Qs9m
9zZNPf5Td6dZE0geM0ZcquWEkCMEmwoLLExmiOruu9MuvlYtQ+fTSSr6r/8NG5A2Q838NjMphcZ+
6TaoQIDMfXsYDGwb65jbqe10sfjJTGUYBdjDCKxKgXjL38BlKm8lt8x9rAwheJtreQo2U35yNiDA
t0HVyzRx6kwHgYKOGekuNy858GljXH7gvGd/Yh75Mm8AXGRJHnvxwXtEWaaHtCeeDD8xeWyFT/2I
b3fCwSPcR9bY2R5gZdrykz/WUE+j/Uh63Z7Y1b2ukyF4b5QFilzcv47RdxJpHDAMf7p/mKTXGfaT
V80E1p34GWU/4RFM23XH0VcO43HvBng9XyfZpwEZg4jdT3oGVhsH/qRKFCqST+X/SRnIigwsshWy
D+12lRoSumdaTCm2kvv4S+h6oJ7CE7XHIewtMJLXjThC+I+dm/6O3Dy9LTb3B0EGvYeegZTXXdrJ
hj1zplU6lVq8PsQYVobJaj8lhzm5qHgpJSl2x0eJM0drq3iXmZnfP9soeeSMPyzPMPY7NPM1FJpk
nT22Vp7yKqoMq74zE9JLLyiaa1pAOeg9VS2JjaZT/Hvoq33opxDfgU4cmLAThiJT5F8Om2mxhFCQ
Zd13gZLvlNfd9T5Y1cVDtsBlQPOtA/qkLJ0XiyzNUcxAQiwtpt0qlHXMJuF2XQa3suPDbaXFoAKv
zj75i8GkSTgQGqmlDn8ExfHKQ1h8TnnCJDZYT6EWyOxjhzL8x+HNl1tZBTpzahVVRx/K1qA5pXvJ
gWmlc4HIF/HtAAS/EZBJdB6GNn4gT45aMS/Jh4q6pdrU2s9Pq0SHN9uqjVdhPc9gDJIrWJfWXxv5
lUMZoPf24BP2df1U5GfPBkLdN2W1oQJXc1cITBfJMb14yJMpSfWURM7MQb36lexB4UfrZtYaIpNg
lPJGPi0bA30s92b6J8bZ9itmUQlTHFCGfTjmFiu1nXGZTMTXpG/F/0w8wHXaTiOt1x+9yujb0pcc
hkaZV0XIY0HMbZ9iLUMMxaGN/gpyZqHnoF+VBwNqJjodoIXlhR02tI9HovAZtKN8/prFMjvlM0Ca
40hcY9CY5UBCO1vrJ9kgJJtFY9BRngXcjSjOG7h54uGVVQ6+CzF7aZ/LMhFKlyNthPj7ZBaljHC8
hLAEqHZzh/G+FQEaiYBuWG2EKJhH1sSWosWH6RfCfwbMYjY8kcF5zkS8RuWXYFY2Cbur0R61XUx8
e1uRHvOvMHJz0MxadASItvyPVO7IWxF3jsev8NQya/KNEHFwbvi9MFFPRIKla7eEJ+b61n4UyVF8
QW4EcPZTH3wJFFC4sZZ1cfAQ1Ex87cUlJPz6/vRAH9depS4QrjzcQFsPPcOam69mC+9fY7As7plO
7/Xnv2muxW0a/IbSiCYXKI4No5q+rc+t3QWpAypIBHYtppvDL8MdRFEt6DH1v/0T7TVh5iJXu4Xy
vhb6/V0zu2jqJajtxFpUcidQJFJXZpG0bCbhjcPV/uyvEBvIvoadGTxBO0duAqdWbOQZ8e2V1k5p
Ex0lcGzC9ndxPDHn4rcqVZRdiaiK8lNjxMzHmYZkBA/2fIziYDksf08L7Wc9xPyQnhyejQK2ti7r
9YirAARxfBl+GeE3AR24cFGFKQUUI5qfWG3aLXV3P4Ii3vWF0jK0hNyyq5Rc1Gd6vxS7M+boxbEF
YPR+UP3uwAKbn3MBVU0gSncerGzgGbzzLeyy0krOcTsWjz+x6jlLVw+Nzcwuj4AsNEBSfO1FWisp
cO/PZSk5KxxzHkWwKBd9c+dxge5zw86yrTKmSm6r7796r22TNQJUMKZaEnURL4FKFq210CHaZ2kB
T8GTxaWojs+dlFlPp7H1PNtrpMJcz0DYgw1waPbZIK2EZDbDttboUE4Pki6QSRuAhegNK2+3x/mH
8NvTwcIO8c4gTpvgvaXIpudzNh311c835+haGFpRyh2dHQJZDeGi1qdUv2Ek8KZkdLAkWAuOcZWx
jKR2wTTGO1d9xVVW1amyXOtTN4vUutXJpzqobjFH+M9EIiuI+nroRhRIz/yOvHagBw9cZ9dX+mW9
+hWx+tzryjHX6XX/jxqBnUDtwjGj0lppYME4QR6YjIkEWFRPIwvNWRcwgFq8WoYwwGwD48KLiK0U
Taudkd2NKfBTKOETJi23sDz4QWVcg5Ju+tfLDQkNz8TF0S5Jt/NH9AZebnGVw9eBXF6XSyIcCt7O
36+Zl2YmtmRfQ1SV7/WEtuhqbUJPyaZL4+Ywb4TuWjUrFBYrAg0b7R0sCX9HlM5moQ/BjrZfGJt0
1RkMfxaWXS+mgemkmHVSQK4IWVRptdZxRbhdySiHWGJAZYh10/DhTCq/0somuaoU0BLHu4AwZpI8
rKlVW3x5sR0y7QHQ+Ih4ds2M7sN18dEUmg7ao60FdqONcNlglX4V2cOh9TfDNEreOh/uO9p6kZp0
n+hyfmeDsTRuBdDoCHnmFe1b0AY7PyYLKpo2SPvtcprS8/oJpKOpmSTkbMfUerVnptZ9WlOS4raf
ro6OUIzCIrgyVrz+SiktX21S7dGau69kZ8ZWbLSvLaVoop6rDq1PxFH6wlM1oPVKj1TmsdIuuJsd
e7bo939ciSIRNzqXS7docB2xTvL7qlLnHJdIah7espp6ggmDpDeQugc+vu0JXddGzxLUnT+2j0Cw
LFVf9law0vVvQGkLkZXvG3Mdjhru6jWV9iN/TDFwlY47BbDG+9RlIoCJBtjmRXPBBKUR/nAdjH1T
CEe+V41yApTBm+jbujItKFDrCe70iVBp/AM2Cx1f/jeMXzSzvatAFXy63fLw1zvm3YP7fH1y1Dzz
F9nU+3P9TY8tNxgSM6V1OZIsKbrLeH3iW2cPmp0Qhpg8LPhDG89UdQCP0TJ7PjOZMH2EOyCg785c
9okDkMMprUydFZXRBEGEFErmfduEh3OJnLxdsNufS1ktlx8iemJQHr54ioVcGrGNV4T3s2wz8xIN
+Cirfvdb149nCIX/G/4xpAxeaUu81RxCo3Ou8T9zMd6vBP1aHmqWLMxmb4ldJV0xdIBsfZXsG+Lk
3cSl5EwFEkN7BVlJk4rYAYkB9w/O1Ntdv4XaLz/7ZvyQdnQ8l2EIwQknVWurijdD1X1455w2u0or
JU7w6EX1vYYpuFvRKMT55arZHAMARJZ7V17nRDhVCytnOc6tLiLxHty8C3tqCy/D/67sJ1dyk7ra
Nn80xcqTzEX9LDrK5/oin9OmrLtDU4mxfpxqGOP32xqDhKUabbE09Ywm6NbPYAQRTFhebLAa2O6P
n7JdCtTbPOzvBaqoaqVqWZUcU9C4t/NP0bwOzhLSDldKB9Oj4eGazYstA1CjofGA+mohrdztlN2R
Ool+KtpKup92yskVTqnQS6ylLLrPLK5bxX26MArgFQHPcvzTiEN/t3SuwM1tX29wxXglxnwJe1Wr
yWSscIluYNSDKc15dYdbgSlcA3vJXx4Kcl4UtyU9npRgS4QvPiho3+ATnbGsjkP8upo5ncpVDq7x
OKIFJCcO+2vGIngKKccelfT45JhIlHMX/8Af8J1IZrIrMhkfpjneDxGsfWcq3MQYtPvGILsyUY6G
LkY2e2PkhsAlC+Vfb8vvPLJAl8Mk7YvELQ635q2By9SbjpRFLeISCu00WGHpCYQBQNwVTIQks7wG
4Gr7EFzAr58+FqXoma8yEWaVWcR27K+0fgpRAwx9gAL1bsZNAU5tNggKg01RvZekZL+zMuGl0a9t
40nmMSSIUauMK59Yj7y+L5WZt+dibEqpwAhZT7fci2KjCB9wGUNm+f4msjzOmr+qhykoKfgjWdDn
f39Nfe4W9G4wAuMsq94+/PQ0ZoLQudRdfYZeB1dvOw1sJdJshdilsZUyM8rNze8sT5gBqQ+pkRE/
97+DoJ3MUbhOJRWfYZFkxbwvfltBlwVF+qTKrvPwWBVRPIWNU5K0Es588SJZ09/TOxHRuNdeO8Yy
WnXevYe+gq9Ju/woujHLeRRSOzaT7jf6kVbxYZjQkfNtqaphJc33LPPaCsPQFKxllF9VKV64u5zl
vvQ00axjuTSnHCcWpR7ewAnNtpJoC4fNoltbyFlWkQ7Jrb0PcW4pvguVPXTMLXnrMQMlpkUy3hVL
sNdIQI/9/EHu4x5Jli0b7uw9jHIalavfdj1/jV1CTbGB6GxezdaGE74w0U5w+AQkPLj4Z554eiOQ
hF1FjGKpSjzWMs57iKU7pjkAI9rnjJIz2dK1ypazRwN81J6uV3gITOfIyDaL23gnvO6HkaPzdu8/
XwaAz6iTYA3gZ7eQo7BuFfVrpv369PsHkonJJ/htVgiLW0mXZ7Rq+pt0AQwfUTMXDYOF8gb33i0v
/b3ALDZuRnV1mdwO4jhvuHbKH6/4/3uPcVsGDmq+lJAJ5uOLzjL9d3Nt8WYMTe8GdUe75Awh5Q94
AgrMTufhASAPYr7W3iYItd8eC0o2VDgjAOUsJa89PyfIkBfwxOFVgbQDmlIrdAA6PA3g1r+MLaHF
gAVnptEsDciFB9ue1Oa/Vzo+tfYrJysTOXluWQNFDRLkoWPYxRbqfdP3vW/YOtI5B3elaBF0AsyJ
cGdS75sAUgzsTBKYlsBYNHVRTAXjFfMrbG0m5u8u3ni4rtwJsi/hoK/8eZ2wCWFQjoAL3/v04PX1
ceBRioZOZhKwZFsqD2/NOpd44crNakRdn14n3D/ANJRGsx3dqR301+dvDSA41iDxQcIh78BO5r5q
tigU0Z0Uiow3Zl16LAF2jbikCl9pXqIL7t6B9Vw9hQut83yXPTh6unD1CJLbUVJJvBJCNfUTDzcH
u+cor9pZOwofx+avzth+MTTsYhnCtNLJIKBXfua47TLAZvl30rPDzaKEWiAOhKfqkhYinJYmAZc3
ewfLohxs53/2dxhCo5iYAE9dPL9OJSZWZIBgaK+9bq+oFB5STG/GKcsuteHB5FcGnOI7hLCyk+bx
UFWhLO5dHvJMjbUCaYUSMMVCNaV77IhPLEELpuZwaBEU1MYD/NZWhECVJxpZtZb7TAfasYERCcUQ
lUdygOU+Cz+4pPoeS1sVskRh+4jsKNSKSlwFmaqG5L85n1MtWgXsdPzFsoZ168eFs7ZmHhrtCi7Q
sky6d4mJhucpN4rSGb3m0znHoR9bR3XxPje2CNMjuUi6VMLxBD6SlKhbg3ABPE+yhjHNwmCRJVPi
PQhkfg8AULgHfs2EcVYpL8LJP3uSesI5hCIxE5413oTgYIf+J6r2H/t/mXlYltHBj0HnDr8Pukwa
oZPFG+tXrwFo3RiT8HcH0MU8Wvq8gUrnyLq9s9ngJaxp3tYEyutx9B5jfMeUHDBPM31A0jhn1IdA
skDyuzrPxscu/fje3mpsj2IA2fhG4NHbICBSucTT1oSjnBzkMyPc3rf1L0prq07wZIkuo6oHuLUu
0+vahJLOod02JY/JUeLbALPhaC5xz7I51oGEKuLeXGso0Re9d+amy/NG7d/Lc9vl7b6KvtR9rwtT
JT9wTS3wQF0h6wbQEeQlGi2ofQol5Wo8VTYrU4+jz2okHMyj/OQCzyE0bZzcEbajqYA7KW5qpvfH
cm+XHNURb+ksUSoslW6fnivAttHuteWoocL6Qkvvyd4NVCZEDVJ0/cbn9krCOc2UPxB71Kl8KJrA
DXkGy6+L4BnO7G8g9x4lDZExL/935Qidilo+/auA+1LEKySluxvCtnkp8+MqetmIEovwHoDKDv65
RI9hqrmtF1CX/nf3Iz9JEJU5atewvv7Ff8v/EuRTe5ByHQIk5cyNribvAceKaGAoRinhL/6DJDrc
XtySGc9Jx5efWdzH8iC/Bix73rf5kCrazdOEgtG9TWdAe17jZXV18QV0+L0Kz8CXAlLcOF066akv
QdAFhdpPXM/DlGJD4c3gBgYjyaR22/tIXoEZIScjyVRe/r6NT4OuNcLIoyYnI2z4YmXSpEve+uja
6Dz1Hm181fewlC0XQuNr/aTwaUl2KaQ5YAv9eyRx6KN/0/Jz0PLa0sNeRpzVGSoDAfAUgS4IXtCm
6BEi0IURgMl22uJjWf3/vl6rpwT767NQylByyQ2galXcg9lBi68ynwrcNVc0d+pDmRccTkOr0ACQ
ErvcKi2ANEQBTnmBG6De/C3cXKgj3meav0YfwWheUYKV6jB7ibjzr2PUdNi+FHT29Birep4QzFaJ
JIlH80pl1Z56gTQI/qDwH4bBxMHQkzjZLpZr+aBexo7i65Ix3aHnnJzIh5SxZYuxqB2wCRfzP2pc
panPGxWCI5TeVmQo06gz1FLIT4nPISjBRa2uRjbDcmn4UaWBwbNmmuDdFjq1C1aX+LbIQhftBmEA
NDRCy50r4jP0o2x2l5UdXWwRxV5REHGVcZ2/rJHw6oxhFQjBcL8/qlikwmQF/Xu47pWIEFN+ZEJF
tJ+JooQpKo+PV0mIjpxuplCo9C7uT7l8JL9tkxhtaeKaffHL2fW+1l0UxyEDVIWshU1jkrGhEVNc
e5HNcmHVkhqPC+0JPleQl56LBL61rB5l8yaswQGCfDkDYSnErDIbY+/8m0ykfZUk/V2qZxCP89GA
NYrCkruZP1UfdGyp2fWnQtbWM02EkYa76s2oAvzBimKU0zpwXZjjr4EwPoukxBx0CA8RHsahQw+d
4PfOrBBVznX+1neR+z1ZweGYmlnXLwSDdaCBHdpfHw1L5Ib/0sP3unpMp9jYNqaeFcs71MWoqs0/
jtslbyCWf7sO5zmz4JO0v1RyEz4Rt5+awAkB9RLVGWUmGrnx1+H7Fra/ZINVjAE1azF2hz7THQTd
UhtMdOJlPGJOXdWDXivcchKunDN+qgM9Xned6ZbBcR+vKNLugLgYCRV39oGFFg+0S489MhIg4b9Q
qFpgS7aLmQfDFkyVws3Cii8TUVgdoqs+966Ukr/Lz5fmw+4VzY9cAbhXTFAyoRdjxfs2r05w5CgY
D8Th5ByswjzB1Y+zbAOsvRdcuh1KGlMXPe0hNTse83v4mNRwLcBUAXdoPQZNm2VenMjhXJMrKXHQ
8iirj31wyOJ+VkfncdbMbxrZG5i6tyI0ANp+OR5rKZ0ROIV2hH4PuczT7YLjDe+8y6j+kKFpMn/n
tSTAOOMqYlJF02GxvbMomJVJLUh9JRvywJ+mhCTULSrvQ9h3OiUHTZ9dM2vXU0jiAGfXnejC77zS
SD9ZTzzd43w/3HJavel0x3DNGtG3PD8lZMD/mtNmyjrtd8quXnU7PCbHP0jn7sxM9e4XYSOs39vJ
CtsABJxnR/JK/uxkNlLCLpNQQp73y4Wza5i1CWR+6cNPzcuZ/jtdS9eF7I6fMN+XOx5i93ei9VcL
pbhgFviaeJlEcX/MJrlMMVLglHHQ4RpfLbRYJWtWem605F3vbE2wEAtU92AKpv+8iCAkXS6JmVau
w0S11mPLwJZGbh2rEsgitdfK7WS8E7tezdDy1rTjoCQ/6qG7MhsTQoHwbwFBc80G0Ld14vX+74/F
B/CyYoWghZMp+XThksCYvHXFtVxAnge1QeVBeZ2wtIEKMgnqi3p4QTmJQNnP261krLKxoPrlvLp4
gEdqaAKPW18nnNzfIfpk+s3+FT0m/62bksOnGUxgOVTkOX3Dl3buIOUN4H8dM66rUN3KAtII/lIK
8upMEhhwUDkHPLsd9nitYBaPy7lYutoQu6twwb/ovqVqgCgUEhG3kXKQKqDgCuO28sPhaSqzzsPL
X44JkqSBkBwoA7j8mAfYR/i4iZ3kn6gRbKDn+P5An+NQHbw/f9iBF6LaxCxOSlWFlc0JIbifsEQn
mIR+J3WJuR/cLijDVeIqkyTvxZMQVF+y4OpZ1tf7FOMbn6QrzpiBoHXBrhvAEsEpeCmvIBujObCs
4AAsb4sgbDwYdCCQAvOFuCyWEIyVb+TJ7ZtE/Pykygbt6k5Cu3m6tVJNjr4HUq3xtOIhB37fp4cQ
LNdrF/XIO8DPE99NIizNPAzTeQ6seGnS4w2eoyZzkH4jwwix94fBYFy8IqomsK4t5tXzxLvxeo4t
OD4yPY6sK3hwz2IYKVzsxmrgG+7vG8iTxnjZutNk+YBDZvNLzbMTa29lLKaybUpw5q9X94lDJ3Is
Qj0al4eReAIqNB/6lWdJBNGJsuGyEJG8fFtR3FB8xFsg3rC/WE302C53jqOmin51L+mCur1ypNsQ
2rMpE7eNxnYa4Rvc4SX2V7YdCBm7vU1BA6um6NvCHTiXi7ZDOMeJfmT4ZvPI5NZDspClM1X/gQAL
cT4jFor9q0iJI9hIT5zf5DXgTvOuZxMIfWpOMJhACqAIi23k8w3oA6RNph1nmonS4sYIKrOy6kJE
jJqOK+Pk2pDlhxW9jSWqEPKlNl1XIv+Tv2OSSgabWZ1rEoK8MXHF6JwfLH69KhhH7LuGF9G/CrM8
/i5WK6yUMH3RMiAnnld8E3LgC4nTxQF7cur0r5XaLZM0TGPHr06JNbBEDfTFD3ftn4Hp2i0WTuLb
AviIVTu2IE9w/6H32ya6fPCTtLatju/qk5L4OvuDplaiqRbTSCBbT9st1Dh62XdfoSZLsBeHrBRM
X+V7tjWghM42HVGTc1A48z8kDH00J1lx9iLzz0NCwBvfQ0NfRIx+qzJY5iUdTZJdx9t50sw5boqV
BM0Yka/7ofB0tYaaayxNJUs0/LXvni9I9B4berXzt1ZCrNt/LMbENtdbbW2vHhayIBquDfiAi/BG
hHf6RCUaDG8gGYZkdUMkzHKFKPPg9gEMNecI+5SqPtuDJaGmldgKqrwr40P2p/8aG/4mqxQOgLIJ
xSzFB5N0uYKr92aeTcBVJGw6VTkj2FdzRtRsqrk6qbCSzZyZesXHvvTCztgm3hdtdjK/SelvdAga
0wq97LlB3OD+2Zqm1Zma+LT2bnEs7RGu5Z/1wSZ/CjxjkwB9Co7J8+QHaAsH+j5Sf8bK4M0LfA1v
HGq2VYfDFq4nQQv1isGlrEWQ6KbxCfw2BsbvNhdSRXJ4GeDclnOsUxhR9gSUl6jcGcaAlb0tGqJA
xF21yg1UWyVluhRdpwleanA8qRXlMex9HdW0uImQ4+gjOQbsvBPLSDqipLecvTeMBjESGBJhZg/R
aTqoMUXpQ3DjEUup7lOotsjiYJiPq3YvrdwcZiGkB7eMYjPiOwzzwTCp78Acd8c8Kvl8ebVs6Obl
5OnAKIBhRoTKFQtej4J+TtLqYCOmj8qoYC/9IQiMkNa3eDlUEv65e4nRPkz7fghNJgEqGhGL+pyc
+5pQ2narrjbKnzZlQZWEVcLBwoBoeiA5Xo/FOBrunbw1MOPLIpFfHGH2Ekqyf+kCLuyRT2zViref
yjP+gmW0BD6ohBjitcTsefwaBFT2T1Wx3kjJ6bmuu2asEuyibG6gzGcHnB+fqmtNSPnFVdfOYVjd
jQ6cE63KuU14rqmdHHq04eCi0BaN3V0EJg/c2otfGM8mhGPiT82OiaWIP9Xxw1ku748yIzveJGJ2
OPFi6hKwFmzs5AjzQ1L3dF23s69JScO+jNx2TaaDFS58yzbzEK7u+/65vqNeCJ2hfOMizWmSfcTu
NnShqKXjImEcfrf8LslnjrqKhbiABxsYysPqRNW09avZzsuElLlJM7Xk00CHPqkIw33VkZBJaFY5
L4YSEfKfJ+FvUH9BEDb0FGzn1ZzaOZD+igvhUHLpnunv83IxORfOVFUGSV2YtcUZM0Znr6rxfvrK
Wip9DBeOBxH2ilfDn90oxUlwlE37F+K2s8zly9n26WuSklgDic0ODoS9Nk214eerdh77ZZ6gX9Vz
7ar1sQiW7Vn6S5/o+KyhGbViv+RfotcoPlx/SgoCc52ivpazsjhAsUsgaK32gzbbux44P3Q5Obib
rKkW2/WE51iyFz85ckedh5TifRihgB2WoEHhtr0NKLcWGtqEHiUXR/k84JkzBa3hPQHo9DuwuSbp
bteA/puAM2bUBcTG3YFc955rPVUyvjkcoXmMnvqd61zqOHmU9sp4UTDqc1JKOryvGpVdvK2XJYRI
SB08jcY024y4FgCZaC42/kpFElee7K5s/2vjT3xF7THY/CdFii9V0y/Q5OXJzIvXcDvJbq9qBxod
2doka5tFtc0LANwcGk7JUq25PMMruE33QaEEcYddLOIcKq0g8XFdYsFHCnMUep3V558llQyKmQqZ
yFOx6SviJGtRqYDvjJJE+z06UPCstP8d8USc93UCvuxW4OJi1qYRSsgd5Vs33vGc3P7k0CbMcJ6J
NLXS4oIy+PTMD7DvLSwRWlG5Gc40SYq+Dmt/57Ph6TdMo3Nh4PpdsFPLQJZRvMhOPqpQCr7E4mEc
5qbnX8m581iJQfgleqCUyvHOUKDylF8qneelypoyZPMDVKRPZV4KTEvfhWRH9+pe2HJHirpWUsWG
2C0LmEla1ZcTYy312uRoOMpNwADjEAyhnMZGKOwZSuGKpWQf8wvLt7m2sDX6ccUr5lzHoAalnL2b
uboSJH4SqwhNKB7t0vcJzL+f3yFJDTxQ0yBaAT1eJYF62AkI/X5T2/lOvoTlkM0Ij0hl4S65VMcT
8eMUO76ZwWvuO/fHReWAVtwU3oiJC9gryOFhC/X30BcQLni2h1pdaOpcUXdHvPSy+MENjcYZfenT
mYRTnPTf77pPNwYSm0vddBQrDEm2eF4pueb07GlqxoWzF1iuZQv97ZC0PANXjM2FS7RnX/BYyjjJ
5RgIs6BKBJqSEqhtJDojfmVYrt/Dbo+6X/CZSjC3SncxKox14j665nojlcETUpOCVEY+WgsrFKe1
eXVNNGEM/0mHLIdLOWHeJXRmMxpfDd4neZNiuMmZbuHjXIv8N9Fli61gA8L2+3YaKI+gxny4NBhD
Kcim0BKoHoQsxQP3ZsuJ+wYl71pCgno1HA/YPwbZBMkd25bfQtUjntplBiwVOYFy0CGEXumLQPf5
0FrHC84GI3UaF8XcSDCqKKd4JOM/DFHR6eRugR+vfqJAJk2xMZg/rCzkMd9MTnOBITBToayw9KYE
yT6a4aBjXFwbYtqmUZ7iX90qEoqP972bbhjhwoGG6GPIKjnUfGnuCvZQ/WGMJ3W9WNRxRXIlV8P2
v4IFN7cDetUqv3yjVCpTq0fxLW7wSLxg1B1Wmilb3LBIR7Hc/yEOWVlYpRdLozaIr7vdgJvuDt9q
uKd7Aw+CF/IAA/7f9GTmhQQ8Oc2lh/CC54kQXsRkfHHLaYBEb1gnAMRKayasVxYnpDMNXnIo+BOH
fhNYqjb6B8TbJnrUXdUbQpLcjP8LsNeG9xVHM6x8h5iAFcpgf4LqqZNx+0Iajfn/YE33C+C2oHKR
wdcMbw9rrbI3VN79rL5zKoMosP2RV2t/+o/mJZmY5LBzwr1kDFewM7dRjiCttnzZJyF6/KW2dcgx
hz25AQcQOKZ7LKqhVFDtjIIenPXIYKqZcbvgIdeJwISBoCT/pfQnoUAtU44kfVP7yEU3Um5NHfBV
YR3pPyUWiEJgK0pJ24DmOMZz4ZRLVGCm/veNL7Tx2Le27qvZtAFIHqAWUReuNN4gO4cyah9cERTU
xY6I+HMcZwcjU2j+1+teKGhr1IAgMAVip1Ya6k4V/0DQo7rM71SkRKQBvEG8jaxPD6rCK/rSbnmo
dRYhRQbEn2qUViAHq1KTtoWvUC15gT8jFbn2KVHe+V7rqkhuNKRcbxszyBGmTuGIbQ7yp1m2bMdD
cgSk0iG8oXh+s8F9gzeV8pUS3FmPkFRJtoBlKakzyC+UJfjYsQ6bHQFK17H5Anizrj1JxeYgSbo1
iCoqmUcpESlBT9R7KdVKs1YKRf2VdvZv+moaxo2k7ZmVC5i6FdnsW8F6esOn9+L5FMpt3TrQgUbN
AyxuRfnccH9ZBzU0YsBpG2M7sh8V/tEt0WQJaB/MadDHjOQJEe8PkBzozIzkgV75lsWf5JDo/NJK
nmH/lDCssenlZ4KYoxvUn5zTWxO25i29WsctLk1j2kEmtdYTO/oSPN6jFpVeUZR48ckTCwJ9+a7f
+QbRB9wqylt7bx2EIxQV3Cp1Mk1OUd3auCy+wRJo/QAt5UFYbUjmD63X87mKk2SPYRXrBWEMQc2p
4i/Lb5A9wSfotKIAkfg8XjoWYkq6jpv3D74SRZo4+YTV3J8fEUd7ybxXueXb7CNwu+5/ubgXtosR
ADWjpBgdL8eQi3bj/Omgaqgia27bL1MwwZ6sAW4FblFc4d4Tj8FfJzhh0Rei+oWoT6WXUTM+CXiT
OdDA7b2SGd2GHqPwtBo0XAfMHxcYuQ/EwdWQG47cvL1iMOrKe62SvrG+TQSoI6PiDCZpaYKusGVR
/ZNzEa2RxGqFFw/aZtTnZf7EvB7v6QJCQeu80LVrHVleHYALoxkP2qNfGHWmkYsxjCmKiiodIiMr
4tHgBWXPSBu6DklLmxf2bCXbRpkLmEbhAdHG4M3K4eeZSvfS8JqJ6ZqQS6y43gd7Yeb/Qx5Xxjt1
813xp5UnhONcpXJsCC436UuWh+EPNulhcF7+vesVonlouBOlpACn5sahgG2DNhzHK5S3d/rGfOG9
7rBEap4BrnVU7pIwwIosf2Urn6chvso3i2Oy6SCEYpetc8G/yI4T+r+EfXd94lhyMYleSF1jb3xT
mV37FV3FsfOZkPExuq6ZEh9SGpc3X5vw9UgddoqarN63MPNbbZAyN+EtoXgsMow4DTbCom66f3VW
fpPnHyJl44HzMqfr6bVEnSIl8OU5FrMtuWlbkjAH6rNM0A/ftZ4E06wjV6zsq+AtKGc+dsUxXJ6K
ix4vvypNBQeExV+gkGmFY9Fl+JbqZahC+m6q5YbsmKN7BRBZ/jp0ybKkP9+LigzFMGUz4NyN8DPg
5SIyai14q45ofDGqXgLi9s/FL5e94K0PTjsYr7aPhTMxRj1WXwONVDPY4IYdgWDlv0NBv1d2SfHk
72RKkn8QmujtfhfUEQyVl68mxXjx8hW7GW/4DLcAE+OAKjHfY+DfVsHRM8RF11xUYJD8rsJ/q9rA
PZ+RNgp0OqNNudO0ABl/IZTu540VzPiv6RNu5V23xcNUvbDIj3IFluRzvOIUWFKZN16/bsW2gW7r
VdzyYeWGX+yivAtitFaxqaQu9U4f9Kk/pKqe7ury5uRy+OvKQqk8KirK1MLEDSTaHqd/+rev6c3q
Gh1vclNJVms0d/hJUCgbNXM+T6vfTTcNY0e4ybMZGpFRfFbPtWLRoqvfFf9Nn4gBm/IhvTxev9cQ
3BRa1sCyoVwrqJC77Br0bp8QTcfAVHm7GsDg1xBJxcWV7MUttHYgKpwR7ojQY+DosaaXUqJOziir
rIwomoaAxj1BihWjR4YFU0uHw6F0Wcwd/zW8mu5qRavFY3JjFfDDAcwa1u30/nPHyBF1QpFmqyUV
UESXMFVzoQgiYzpbTRglIXY/hJufApIOmefl24kZma8NKXbW14iKNBBnMA7Y14RjTz8Q5MYJ0911
UdvvYlnOJ8iiq/QNtyMSL27faIDbjr/oGli6RcfzPhvNBG5JEEeO2RMLuT6KSmSDJ99i2Db5+FmR
v7GaiY62Ao3o+6HJ84U6KPtjDqg42pEvUeOIcRTe4trK3xgsBD2vR8P+zQtRIH8kAYiijO4O1+TZ
OFimze955Hn45HzdTRkdaqBSRCX6V1eVi0/n1csNlBW/rpbmVmBJKLpzIIKcDSX22yIDHg7lqAfL
klegnaBfZBRDWq+W/blR6VDf/Agha47GWF7BDiFTxSdStjUkuUSG02Dy9UCbiMkdEV9+yGMwceoy
/Y5+a4iy9MpIshNuYZwBlkEk0mNbtY/lPWVhMOoKdmxl5JnulGZwmif5kv/pdbqI+gIfbu1eQ/0j
xMscywZxxnIqaFo0RNSZa727126w4MVgHvGMUUW5kf/VgFcYyuEAe/Qz6VXAyKijaLcJsr3KJIhN
yEjZtLO90VaBPwQwzJLGN8VuUYkocBwKR0GmJigBDQjNJv0sRBDvSSEL4O8Ra2lGuVZKGm8k/6+Y
osLcYi7O/4VwrOszkoM8X+vXPX3ZGK63+03gsXT9ce6dy/3bmgeyw+FrzUyc/7iywlFNdWNG91if
sKzceP3qgR570bLZZqe3U7QsY83Ji/K3mVgKcAduaWqgsQFMmG25L02rJYlzvzItkmomuSt7Kyo3
9lEG4SjiPNwcDSSvZKHvS5S0g1PhMrDilWVt26JE3jzzAlh+nSRfHClZv1t5REvCH4r3hg2PqFri
Znv/ltCLfMeS+XwHUmXmOz45w12mfjdow13S2+XeA0ejnfvvhDICM7lZFFcM3X4UnBlJrb+1fs0v
Rul2Q9y8cfJGXdIlHmhF+gWplj6RgU+sm7nECUejeIcmk13zv3fECvr9cSbVDZ7vNPVG9hCWrm/9
lgQ2S+k3Woi6I+jXvAZidXj1aHgvVzxsYD1q15zbp9mP/mNIy8M7QH5KnIQiW0f338XLWgvNKj+l
rXFCGG+ymVFTSEKRWdFEJEeUhRDtfSETZrPq9lrypwg33q58rEeNg5+SMxTJr0VjS5a8/XLjCKxB
3QLyPW8Ga5fb+EWh5mzOXZFdUogLNTlrc9LN0RkW46LHxgYeT5Hwz0NwT02v/TtP/DsdjMQTbS1y
dLTciPM1n+/8UJq8omKX6FL/aDcTVfEw6d/z1rRHRmd5P3V7KQAPGUn0laYLMespTUYI9X6R0n8u
3UQZuZ2vSTnCUj4PHyRoRPqc1pQOTlytOVT2aLi8w1pJTIR8UPNvYD7poQoECos1GX38+jGErksG
mlso3mo37mlrU7QOUcvHxIoonO/hHNBp2MO5JuINetq1WYdMCkq5cmB3ZyPTOfFuo+zrFQXSdVzT
OomK5VvSzqsxF5tZHja6/W9g+Mh63hWK8zCyB6RNoBI6vfjoWMYToECReCJvUmbIilgIAMqY6yao
JTJwOQQ73snFpqBdo+erUzark5obLwf6tUwojOvg0U3ufyqpdtDSpELhZEa7sOuKVM7j82Y4BLQQ
MrZDR9e4FV6hbClYFQrZ6fs7/BIY/N07XeNZorrqKyjmnDP6iV0W3UAh4es6dvcooKYXZsRCYoRT
AgWq1UnCWWJEs6zgyb+MGrn0pcs+B90H3yR2r64Siqhfv4fI5ZXVt1sEouQnqKlv+X19hV9vTZuc
pePA/VqGUkieN/YcSxhmRQMxUle+G06pt+NNKy32XZXGCVHZdl1JGd/Ts9bTDEv/x6w/B9lxjV2y
YpiJW6PnhG9csbBI3pQ6jc46G24rsG2qw2jaTPqsU4IIpuJqPyYxW7xAYZMsJNcUGnYPmMuyrCrt
YYMAAVk8FNRvOPILWqBUU5goqrV7+6upj+1m9qzv2voNbmGKrsaGEzEtF5WU24Rs9XAt6uCgp0NG
SOHMXqo0wiueRDiGgdaF+4hDO4Uh2PyVa00tF793Z7+V8M5RE635NeaLZpVhSBOVqyMbay0XWhxl
/PIjJBwAheKTn+cCdTL5gJdVRb1Y6wJWvJF4FGHAufeSxUOBJucuh+QxUflUr/zUKH37y2HH+NZR
K1ATyIbkgZpJzHm68QkVZXMTNmMHcA5EvFzf0n3IuR2AmF6Lw03wBJzjMS58szKW3EPLOdUXKOo0
yAznW+i26wvYpxTzyJwNfi9wX8PnXbLs27O9DLr4FhWNXA3xLO+1VTTE68VMQq6v4cQ0Z4aWvnVa
Wvir4GL/omf6yIYZAKVGIJtj1QrI4Kv9vz+MzAuyBqhUAVR6ihA+E6bjJnetMn19Jbuykwust+zK
B0dQ5EtFXeuYa4ezVswfMgf/+mxCsUW3NgstyYruToeTDI8qQfckClfyyr+4lhq9yr6dknaqM+U6
DxAyws07URo46Gq24o0M8JQI20T7LV9Ka6XPLAVoXZx1RieFmmD+B0SqHPDIyVXwnCqA+vqS4UuX
lY1JuchnO8JHq2M28oCNUZMMEb8Cv5+4TRo9EXlmeaBUCAtpZPzmHOIzbmFeRmU32h1wraL/ZiGE
WSMic2TVcxSENFEqnYvfL3RNAoPKFLTCFuZcm92WNZRrc3SUO3/ftOK4gfj/C/DL6U8GcJIhyEUv
6QNEKQJQ6oKNUTm0/cSHgCbdfDSrUCsgZVGuOF2d76g7n6pdq0Rk2IWES9FUCjcdCsQlh7bktNFd
ZBz33C8GNVGkL99zoLPfCMzX9XeTYuS61m185ymQ2RJeMHFsVKacy+yJfx4VQoWDgTQkT39tmXdd
LiZwvC1m62r82pHtFXqdBYVmlBDflin28O0lkcZbwKDm9IB0OjCD6MyyxRTA+HnjbxKf2lHa2OpG
U13ohSkV3lQS1pjCwNO+eD1qTBryPagtdOaL+0t5p104+d36l0D5/tQmeeezFrGkEx8gO1CaNUGA
buZi47cUgfBwTg9rav9BXsTIfYnUQVgti/V45IuOANiVFd+LKbpjiA96MF80QIJdTPw9cr9pdjsN
w0Hf94C9RH/WPweuUK7Nies5ZkrInmEiIkW87CKhc5a+DHLMutqn+KOfQp/9ysYPAyKRto6fXjqP
5EI30ROAzgEv0ludMAiTiK5ex+VMS6SjyWnn0+jQBWXqAohixWnxGIFUA79kUsmQGLs+4np7Ex5Q
AAkZbH6Iz2zVIChDeqDWjdsA1aaUtykUAp5X68DRB9qhvJS7m3TjiINHR+c3teZ0Ct1Zd53k6m1n
NDxv0VkweklblmZYoGoFhnMyHgtVk9Hq81XFRJMqV1NZH4rpwTH/WK1Xk0CSmcSHXZpEpMVnELu/
PlBZK1/YFHQ8uhhU0+1iKExSaC8Lm+d5gaMl6Ap6XW5kEykwGF/dTuaY4/0/784EoF8qkwraWwtm
WrtxAOxPRb5NAEjuwN0jLS04ozA03QYH+zLBmEDgehzseNnPIgnhMd7i3gNOu0JRQSYjRmy6mH8v
SHWvwuANfoiVrfUjb1HlkPHqkzT0QgXBK6QVn/X8DJWHEBeIiHEYZBZ8IH9TGPrQHzh0Wo6IFioK
yezVG1srpW5elE0B7RRD78PYydSkUi/Nmk20sAu/wJZ4GbFnRRDiepBCivqI++wEXE9TwbLRI1+4
DhaJUqSwC8BF/IbgeekMNPOhtXzzPUlpoTKYD99cZLP20qq53e7sVmtr3FZNwvV2K9eM/dz/0oV3
h34smANqJ4j4yTf0lj0YdfrRknu8yF6bdyDS8yeZwYkvSB7DYjUVTe+fQ4K0vhm7Po32/AFBo5am
cPivFRBeuAgDQByY5ErnHiZu91cJdYjLGteu9Z27o4f8qUlu5E/fZOJ4c0+3V7qVgRNZD+hMzpXt
EvKSLpQFEagRbMNYxE1WM2Nu/YU1XHQwRMm5gTYzuB3vKDJaJOJ+681q6yWlTvjAuXES1UR3gf8P
krruSW6hdzOojuDw97H++hSVw+x0aQvc8QdU/6WYVGb1D1D1Dag4B2s0PXby0b7esldAXlwcyBjY
Yf0g+vngXNrQV712Mp+RKF4gcFAZP3dVT7JxbHr6nJqnyFOwIw8Hb+uwxg67hOu6pu3hvz8UN041
yG1VNj9BkQwEO/pj/Qv/JgkErq2kslD/Ao2HKBqRi8Zybt6IrS1d9uFlz6EWwaMV87M1cGU8Scit
gIqhLLmzfTdPw96jBoOzV8LgIMqmTBNoW+Qj7/JPFswyXum4HsXmVW17P7PmVL6kR4z1iB32flks
IBpccDcxamQk+rp0pUza7rrRBgzjmyCsNUNTx3jvS0QV34+5q1aKVrDAydHlhUdFKh90HYba0WhO
pDiQEUMHSyrKgbmyvMWooN79H6hqu8VkngKovyWjs6yTwHt2eBtXTXi+MEi1FSAvQSKnQSStJq/F
OhM41XJv5ti0apV2g99SHeRzIcq8VTyjTYoAu0LCaTxFHsS7i+aVa7Q1UNT4oTleooutuIWL7aXH
xtQGk8zf9YiUcVxrAl6fnZyR/5e4t+NilmKHVkk6x2G6ZJkkzCJ1HUt1wvfVpPFT9/fgu9ws2+Qv
+gNoeTr09iJP+b8q4v2lo/IXOVyfHYGdASLpby4pDbYaw7XEFKPyHhnHbPXRms+A9mmCv9bXO7Jw
kqG+TLDqiV4rv1VeqzYN8WSaRXnd2uM0W5KF7SMhdT9Td42lUehJDUMm2+K9CgI0ywwRgQkp04PH
Zm3wSHZLvoA7VpdIcIzOSb4bhd+y0LvS1wP5Wm1vj1Di6hHkOrQx4GGuL/uw25zhZyE5mtCJe035
dZMlJ0tsCHyYAMWEjzoU1SUuByf0SmQIv55BPMbWQse6o2n1ng/p5bKmTdRFmXPRZwHOaASGLnPe
AJ8arKsBFk3bfcqOyVS6iq6F5pY6gS7nB74Y5PLrJWBTQIO1X8o4wWap4zdMceNCvH/eG3jj3wLB
TZ3XG3/hnr5kVhxnrzzPTZtYlDff7GOeoiAaqPvRFlZTASD/I0LZvttzjIb5o6cjajvLngCTPiiL
xZSjSYi2a0wf0FVDWS2lIVNI6VZ/dsHvWcG+Ig3TJ0JrsPoQeYILkTwwqgNP+UaN4n5HycLUHUtf
CPvOjhRUOqvlrsZA7RAEwtxdpBKxN2g9o/81WGxVQWGsS11m4x2OOTNDb5IayDcB0VQ0bAiGYl7A
UmlscRWNWI/sRmY1iKZm8eORlIZ7ykwz7wV40aEr40FwFFvIoDPgXvbmRuy3mxoh6QyruKORNzS4
+QC1+x8HojHHAN1cN6Doi7hFa8CnbS4ZIDEKeRp0iIvaneM6UWx1jAqyZ0uWonvEXUqvZpXxfqKg
fgoJ0PsqJRi1/dnA1Y1fM7aYAQ2l/0xPWAJLI5UpCzC8jTXfBTwpFilRfXYQOCPOhyowqEkY/dSC
702rEr0j7nKJSiVy0mnn2UlvTzgqGWaXdEhyopwXQRtzz/uBWrifj3qnzDikbcZ06QiXyKRSqZ8T
qGGEQwQGuIW3Ey5vJfthrV/mI5B68YNykTamHbKvY7JAlAcDN00RaEcL/+dg328AmHiKsuJ4/DIo
M1Zbj1UxoUyLzpABdTNnBuvWe1KbK+9E5qpZS5mTSZn7N0ebG1Tb14TBxqB5L6Kbu0c2Rqpd8OxX
sn0g8SQ23hfPMMGdtvYQxTM7Ye42a8p+qifN1zsSnphS2IomyDJYyfkvns5dCOE2YBUrykIaL3xP
O93XNR0j7gwWOcniAdLMkL/Sjgpsa4zD+IG3z3rkVaX/SMHEk86S6XH3UcCi/tkNd8T0JAutCSB2
Q3RW2TvS8/Aj6MCStyVVgvhWVOV87FnNcuVWQ8HKxI8dlLR8CyASKLEMLh2LDIv19kbLz7pbI18/
jR4EViKmE+VRfCAM3uFZQSa/QTbwVvtKq/3hvuEE85kdxeab+r4ajZ3kTBFX2Bx/s/nyVk3yW568
rUnnHrgJQfBElgCKgO3/xNraOB1ZFL67uP1UcoRR70BV3W4HKr7nB81hpX5r8qpjuPgtMGOLKl5s
N7yawusxNLKOe5QvTfcNWc/oS/NP6gD/x5vBQ/Zanh4P3qemG85TbMPKV5yQjKnftkALdThnJe2V
1FxT+O81lcSp4LRsVH/bOCOeKuNCz1JUzeW2Uo7xtbLUDoVK3SEGiHLOalgc4oxInPdGYWsjRfiS
xHEKUniMGIziFWOUaYlMhukrl6UfeI/livpzfZ8Vi9nw8wxAo+JMiWD1P+WXzchyycQ1RpfGS7Br
aYeVYQRcGPdPujd31hEu8IacSDDBuBYTILHw/OrpVzLIvR6X3p29FudcVVCHDL/mQpDc+fr9qpAF
PN26PQDX1jbjHQA6EwRqy8knpvmyG4ZjlgfjeutEK15K/yUp1BHfI4RxMVM2yUd8BmKfRg8lDldb
OAtXfkjG6z0Wbkr8wgHz7z9xv233yY4G/h6yewHpX2A/n2S2PIBq5x/PqeCLAIx6rDZZc3RJcJZE
/VDMnHVj0xzaEOEN+Iqw2agkEcZtW88Sth12VS8TD0p+YTEX/QgpsgzIY5U5Fiil8vIMOD5xbvy9
eBgxdNRuOyjrZf27MDeLvr5xqOwnmqWCha3Kl+sAZSAeevs6ztDfgZaT373RIK7QkJhcqPkIEGG2
hefDlfruW1TGLIiGdmJDtc9/7Esad9Pg2JeQfqO0Upi2UnCh9tPFsI214m0Ofj4cBh+dVFHXfUfR
ZJ7MRZDl9R/KUkb3O9PVkgsVP0xnwYSTYRfHwRYDKsdCyUO+Sci1a0O6mPsNF/WwdMRRJQEeZmq2
+pfu4rNvUNrV+FzmdH06Q2OsR96Jotdd+RBCOHcQ3v60cqfvC3nARGFjFlvWD0wPw7GeWdlZj2PQ
K+lpkuFZ4hRJzmSzT85+ntj5zLzQoV6D/Dt5iUdc0/3sBVe+n6gdFRtubpsWi+dU8ltuhsVa6kz3
g8WQ+Qs1B0/ZvW64ZKzHFFLe2Zm066kviAyW/KPZcxyDEOFz8yLB+D0eQDQoJL/PMVAxFHUywFqU
/t7UFJuE6DcP/NXsnCz14XU7MYPOc7yN3ZF6g1A/BMs3ptYiQD2iZh+GxVNIw4fdhgF5EVXHw9ht
DTWk6vEppTL/Nu4nXjuwHjUn8VIjPwmtnkZ69TUtXKR3erNXB7fWr4+BWDnvB0o/k/QWFwKUTyV7
xH7rEKktMLTmtfdGyTXYswPKijEQIqo94SqrQx4KV+9nigmSUUckkHcCg5CPYnvo40MBmuEDta0C
QDRlmNnIFdVdUdme0dOerlK/jVP3/qUH16zjLhTJK72IhK/W5SCjw1I8aeWZeaZekoTfV8Gf3Nqg
ElBVGGz3Kb6p/F0hu841qs9pB4E0nvr5c7Ch+0Gu7FiXBmaSoLZbFS11/8V1CkODeTDPXC7MvHBE
jZiVbKmkCgmBTvrDCHGqLUZ1I7C9FnVbLC1Ogb+gcDevWG66vSBg5DQFabjv/5QpLPOchjlNe877
R0k2cCf7Urt7vxgjj3SK20OcIx/Xon35hlPr9raAlil4VgnKKQZ3JP8nx38tmjXYaHL6dR5GYo5t
BmejZpjSSvj3bSY+pO0/BEu+6fs5M6MH2Ri3t3oDme84X+he3EG+wZWQayqtdIrbKFg+Z2SGDV7h
aewgVHEiLr797CWPmfKgjx1YUbydLN8F8++YxuxIeM1IPg5+eg3pZpwD+VgVZApu0NsjrfNuOV97
MicsI5/v7nFsTBwfqyeWEtky8bLJxiDnKoVNFaC3quBtG/lmXiJG+bxRy05qFpf69x5uvXUSYfcP
FWmPQwoPifgHeD5Yk4RcIB173kLLl6xnduWOY2KunkY/9XKidLLkf1dcLy9uuFSRwSN9HzFHKgl+
kmcb68SWMhJ4rxU/RPRyIpe8p0uXlUORQqGPGFBnuaTyHsU/po8rrY5mV+EyhgYDAog4IT1q8kqg
+y6JE2UUQxhYYT/DNyNlB+ZTAicF+I6Y6Z/q/HjXZugBpowgjPbMYPpjgCsqqGBcT6d4zU5hZgAl
0mUY/SqwO75zDPIygGzyKZ7XAiv27o2XUtawjl9reNPmfW54FfY29zD+aRE4itNP2gTX7YO9NncV
OMLWn4v+/C7u/1LUKWPneEiE4hYFtRUQfTmYpZYE+NUwNRSoAuFlhxk8qndo0zT1p+DIB+neN2w0
n/wTkXnrRQsBU9ZWvHQlKn7NCJrQuFzI6jJkE9kHRmjIw5EtmSY5eGHTMoYz6EPvzcohHEac2OX/
YHhp+fmeIrJ07ckrlu5wRh2PX5nLkkUZDyTICLxC/wmxHqpxmsKzpoX0/pmmVmENVUsADvt1PaLs
4rNpnUDBvp3ZqUsNhNso0LIcOqM8tj+rVJ012EdxDjlb9aK9x+DWRYlfK6rq6yRNllPGSP/rtV5T
OdcehCbd9q4UnS1F3fK62tzlX8HgDHOUX+CmgRnz2VcLcJCAmcNAdaLfr3DrgUloWcHD/q/QShTK
VGkuRkS0HfBMAmhwLrvuMpo5PE4g25z0/6f/fcGsMvUldqURNWNUJpijYEqYP7Egsd1p99HoqdKK
HuajPGnmcgprZURIleC18jATMTX2qHUzT0SOG1zGMaqrgc4qGCAS2QFpFDKATlATFzcaZCWwC/K3
erzkMZAWW6y5kLgSmxhdrCFe9i7wt9/rK0TYtgrGakDNcfst+Awr4WkWcJlDCm4909aFiqw9mlnR
KOkNusRetdy/2hudErMj8J7l+UBuqmMQHYy8lnaszoIHSrsRqesAWFSxQYOKmQ7b6XraYiaUNKeh
+xlHiLtBRrkiHycS9h4Wdah4OfM6w8MGDdJC2Jx0LdEF6xjmv0QaKZUKRaHt6nIpoHCcTlNPQ09n
aIbIvOtZfXKTV/Joga25ws2M4riQPKVQv6rLJluWTEQKZpsXej9mn92+hv6525uO2jvn6+i5Qi03
ZMfafoSl9Vz/ppZwA+lwTFOrGfMXdJVCunFoPc6/uLw56IXx2RKOUUGKyk7QZ4QOH1vrE/xFAoUn
KUYyhuHnn6/siQOQSMgIzpt/o2sMdCi99IjwZYE59NTqJR62oJHfTqQGN8oRsFl4rMD1tWXW/yt4
VDIDPZCYWuA6Occ9wU5YRULgOISjC5fFgJsnAKEG6L6FhOXN188ssQFfHJCqutetZKygK70eSES5
bL/ephlP87xjg6uCVLeTUJvpih3rRNQnBDyVCKa9z78Z5lsJeWnmVFfBDXvl303qEiS13OzYed1m
xaNA+cb9W84mXhUV5jZkbZqZHD6x1ACBCQsHeC9lAD8wZcmRufxw7CbTT9BFT+YvdQfbGZhwXKcA
8qr6/ojiIsZY/y+xz0Ggb/Uyr0zoOuCientBuGV5otjwhHNXImOwH0PDFRe+TG27+r5aIhBwDm6Z
zRzmJ83lw3YYFCL6S5RPakFWC2VZBDvyP4RwwNQMS1Wr3DG8ogq8oKHAY7TlsmxmsB+B4XfuY+Cc
WsDGpYwFETMtAR1uBm900QtlXJYsaED0PBMtfxqs9UJq2gvd82VQGGKyRYasjONaH7Vy65T4NYar
0hvBp9ysOpRqO251qgw1qRxU4pHphSRvCIv0YCgORmA6FejaTKvotDm+I8vk+jTatpV0SqJXqDgB
cSjCDhrFhOY9uhLpED7DGpMDSBZshbi41Q0FE5bauUgKxqhPd0Vm8BJkKvtz1U+cZNydrczI+uW+
dKxUdP+8j3mUc12kcU0JCEsIY929jagSlk+duOxK9QlRmw64R8RRQug+LHuf+9RgIwajU9wdu23g
e5G4mRONN/VgVUZRBzKN5qYmDPeTuMe4VGYs2Uhfa5NdiAz48snhVeZTW4KBq3zKyUU5bQBnfc5J
yf+4ovG0qei1e6MAUaK8I7JLksJLVfXc/Ht5ETRoeT/5UEERNKo1tB8MQRkQPVU7NEi+Wpk7hvQQ
fk3xYSJPwb+43edQ7J2oecI5Z92v8AUbe+geaXCZj3RC0w1dL/FRiO0h1ukpW/YS13i9weN+dmFL
DL7OFxtdwCWwob6WkoN7h+oL2gJTgwChvVbNdlktHt1etvGzXQfYjCWgl4zByT7X080Bocc4gpV5
VRNnFiIniWD6rfpapGH4LqWQpMGFr6JFwZBNjuS/zY3nw7KFrq3p4L9oKjsknl9xrzmZs87CV798
McphvrpfFwOozBG0Krwq7VRLEIPWp/fqFmGcLECXthTfQM+vHDee+Uy4oVoAE8btucEXSks9n+4f
1wXEelAh6ndoptQxhl3q1jDDAuH4RVKk8/+TS66aV84Bprf6QXqPrA49uF8iAbHJlJ7J/lLL6RSP
BF30FYK2SNrkmgCGz+LMuxa34/Chq7xiGJ3LZ1kkRWjjBt1uOwSkbh0WLQIGWK2dkSRBFunQw2da
6YCjJA80TB1BlOrT0n4CSrdfpccQYIyOPcvtamkOVpbPg4DZutklJLY+bKhDZzIWA+wJxq4jXPbn
vTJ06xqT5PFTlM49i1L1LAyRJDL7fV530LyiDwkm4f/VCFgMvtkYlJG6idtu16flHz6kiVcgK1UD
xYmvI5JHW+YiaiSLNeataA66PhzDHhMAiqfZETgPlUnhEYrCtcEvISS34EdUvsiPHS8idthb9qu/
8Bn2fySBGNWZoSbYwOmd5Dzx6jcN0BaDzuK8dEN75S0/8l8YghxmK0RZPaX4+qbdZQ+hx6y3XJcM
YnuQE4KEtkU5PZ34FM83wnYEchZeXtaQmbFlAjKB+DJzTGjId0+BEYK6DIO/tN42wqo1icPDQ25P
pfxI/oCp6kJtxSsX8X00WOfcXpSwrL0jtclAKyxXK6Oix9Qam0DkXQeTDnYaEEtyfmvQFCI7hqJ6
HJG+obrcP74jZfxt1RL762+08/z/e0RcbRoyfmbsvhi9j4V8Uwidci+1EMd56XnZn9sJ6YmzQN9A
2PCeBUI8YxPmabiRhvWQfS6wS02E31/vRfkl/HMaXHPFJemSZ/4qGWt59GcgmxUrM83DkC1h6HJc
JwCJL0AwKxIi8cdKp/0NMmkjeG7WjkgPG9Dh1dsJYGNI4+unc9fmsTB6yH0x2kq+0GfRKhw3SCST
jNUoj/MtDoPCrTL9esTeDcWwxlYT+kUy+rgdE7dtzREgSDU+qd9jGUwMEW7AwItAYD5QQmy0ltCW
+GYqhFj2mCRW0Ve2c/k2dLNgd4R2uIIN8nzcoQI7LYGubj9bpPUfkEB6IVE7TJCMTswidJSbF5O+
RL8ARC48EN6J9EK6rKAeWfbSOX7WMyphH3PFwH8net53YjFmKl3favILpk5F9oIWrCSxHKjusUtD
0yBpxNkTkGzDmYRtCIJxDB2pQYK0piWzkM+DQ8PGnTgpPIHx4PErFHpShu/ax2tYCRZADfenKmtb
2DOlbinns/MGlWg6fz4ZkO3PilD7iKMiGBWHmBXaUe7ihJqszSxzzo1bwcd7hFlytaDoQSrOLCZk
2yN6L1QPauxWVBPfyBJo7P037zwE+0GSJNKhDDkS2WtyPkD7cvppGpUAXlJTrusKhZZ6CaU8/cwt
OvX/ugWYg6cm977DJhsHpWlGHt4NZmVDgDa6hvd1W2ZiWD0gVhLWlUswWho31RapFG24bjYFhnSs
cpu2UGDWkwKCRiCxPP2lrJELu3e5lORpXzmXHEFWCqsp1gO0f28W/dM6kWPIkfqLL6n+GO0Wyi+K
3OucV527tl5AjUJdprOGhgLGDNzxBDxB1O1kvnoAWgnzVTaLwBplZskCeLTWeXDj7u1Ysc0CZWq1
eS46Hlu0PmYa0qPV2oscdz2XNwKp9MH8H+jlHyLjwTqTe3lX2kPXMqiAsDFk0oDle8tjde7YPwwv
LUhROOA5AiojuKi4lSADqBr8NnkBT6y21deIcTNArLEI4/tcfITXnwmA+tBbYWFIlSOFubhbQ0Rx
a3hOqRNEWMvXNwuN+lsfY6QOkPYkH9D0l9DR3RFGeVFvLBiKKvAgvvtotcc+UilWp4BQ5X57pG+K
x3YGLt2qhNCknVZCk1j17I4aMbt4vM4vRSFGLRr4iHgmhjbROHRMvX1BWCuMwlQ/+xhACp4+ik7T
WM2sao5hJogd9BLPcdwI0xXY0csJ4xOXgeiw1dqdvIc6v9e8srvGPnVSL1d8dj1ndKe7ypFiIDbP
BArwIShApuVAVU3rt5hwt6gHmmWU35VRMqJZSUKn2J/xnCZzA+3RRndE36MqU1NPX7HcZiqfE4kr
bbZbYRyrURWDxRfa+rYDl9AT3Bm5djrtlsbOe0XAv8Gzn+OXePqraD0EINp5OA3hP7mnQtvhVNZR
cviiJZwmerwFZ6LWXrfukmvMxo8dnF65S4Cm4PTaNDGkAWx6XAoKGPcIyVmfSJLeGmRK9DW8PAxy
duCGdZ/tyukzWI3wso7J+8FjPFMSN0tuyRVd/WkQZqL57lj3nzRg57idTG8zxSXRA0C39Q8+XcB6
pvckzny7JTGafScbAtmRavucU0cuVq3GpxyXnbp0rcqF7Zn1kWhk0H0Ecpz26smPn5fSJtuq0GYE
k1Uqa/hRIRiHzKxjsnCINqDmRyUMP+jsXCohlBOpfXTC5F/y4uJ4zh3cr/Ww9G23SePxZ+76FXXj
h9dG9Dsh8b/QedhIs1l9STXS+cjz05PdpcCCYKdN9FcjHhtvIE93TgHGeBqfyFqnyJ3oHO+cnFho
hJyPQqPPg2sqIKx97A1lX0qZM6/8fK5b/hgROwOJvpq/A8Z/IYxfi8dPND1U6K0vIei+l6eWe7vd
mryg2aeolSdkSRSnFD7KoEann3WyEqLNxbwrWYIaxOYmoJhd0hZ9z4j6V4XEXxr2mo179k+26ltl
KBuI0md6ZRrJIOejPmUi5wwXsLGU9ieIpk8Ir3rYrq2rgsWTTFvJUDHFEZp2N6lIoQK1PWHRrKq0
wn5zo863YyLN1n5L9ZOfkh/MTwWNdQoPBM/CVSpI0wJe2kmaoma1QGyEyMaW+GpNe0O6dbtDC0E4
V15Na4gQWZUyAJ0NICBRanph+lRGWjcPC3PfAFKSLjHP03KoD0ShrALc5URJOfaKN5DNpcFRihiZ
0cUi4RwoQudIuBlWcrJK4hCrQF20QPABoqLY1nVW5SBDaFu51wrscyEUH4vdPE6vxMzAU8e28zD+
zUfh5UazKF5giVfEdQF94R3V2ZYgB1BPT4Wr1oI53rOquL938Pytpjk7gLMpgLcqU/kHrhCXacF9
IfxAVn3f1HgG6vp2lVWzQlbvPF9YcuyWWT57wFiNKyaNAdPgwzhwW+/Il227bTho1NeMMPnfQHNB
pKWy5iooUHTo3Y1Ggi9EVT2fVtmLVYOtmXW4srjcsqz/qlBYSGD/a7ZyO5oya4E/e9gShrbPap2Z
WQOcRyojrtNXNAhMCjK981W6ZnGSFqFhyyGa097uTkr9kTd7Xoz0zGHFV7LglqewImztTlJ4Ecjs
65JxfFBwwBWtGz4UdvJ0+3u2HdQSWdI+XTMEgnIygZZG80Ak9I4Odm1Etb4uEhxllazYOro6yfk9
yUTqRQRYUKImu7KAgUrldomDUqlqXBAklnz2lpDtJbP4nYQ7AbLgw9MWWWg83NVGrIiKBF1HcFAU
HJYbUscsNiFay6ynfO3c84Rqg8CZorTKP8NV96ZB8iQaKD7Nh2gfg+8mQUxNgpz5vGQLLXRg+jG0
pcjCaJf4x8px/XWafxCBEBOcIbYP+f3JkncIo32ej+d1gHDHN1H0/19t6dWpcg45G3Weh2MdPeBg
0/EnGOI4jA45rbuBgQDcUdO2JQPOXPstiipasLFevhorZ9wQQcfmdla0w8Zl/tMfL/jclaFyA6yn
fpMMFpPp8LVAIeGgXL/53miETx8mXk0vc9gMMoWZPheY36oyqYcfKJPieIZXpUEgYAbNdeQ5hlY8
Jyk5eE15xndUuB2zRBpa8AP3bxoU41/TuOoACnBYyDPEJ/mCdyOtvdDxsOWNlp05jEX1DFb2xXrY
e8R3eGTqAfLz75ymI0IDL1zK+zfgi6oMoqa0HsZZnJBhMjGsPCxUUvkQE4WXL/MsOZt13G3jtejS
1REbILepSzPyI0ODhBYc5EqxAkUHhFq+p3aqsrANyQN4ksi4XrLltys70EdpFk642APTTfvaglC4
RUtcO5IalpS6zcPpGIrb2e5XdM1ulGGFN24Z6uZS7HruH2N5sLPy5zAEq3aH/5tBiVMdbJHbVUn8
xULWpm0Lg8q4bfLtZLdJ7THhfu55MCOs7b3bJ7P6lGkMuviwO5q98JWgt9j64A/7r5+tyXG/oi0S
lo80HTCg61pTHT8xNYsHZ7PAHO4+TTKGYkdXnLMGSa0rcsaOnXQzu6CGdzm9RdMjtz7Lkr3zqCVk
X3cF/MDY0U+UO863PNfFxE6PmILP7bZq3BEQcYEn5CueBvtAVncaq1EsUyvFUCdDMaS1jXQlTWNw
LSzXaUrstmuea1uwf4cwxZ+0tLncwthUwMjwfCcikakI0qfnGvBw4PX3Zoin1+CdOMksEaxVSWVb
K/9SmGUlDcqUuLhlOnW1odioio/KmXs7eTRjo712ySdxVienbA233oBoyqaGP+wzjON2Af8cdTEp
/Oaz1Td20HGD/f46nFPjfeBzcNhG9vNtxnOiONczd/Q1jrjwMxAKaCtLfMnNGdc/JN/lLr0jYmpv
dryucvdYCT/7Y/bdu3FJoHphaLDwi376yEH1F8D3FujQXUnllmQiMCp8/RCq5NIfVldY63pxpz9u
NpKnD88QitRUUI+Gc40PhRUSgq5eHjcviiGv4ANMo7wPH+Dm1MSSAUJ89dQK9mCUbNJq8gee2URG
vtAuX1qPNqL+0lr9lTtM4ChAXLn/75yvWE8lrhHI/BTbZsUQM3Si4mSoAqqUux0RBePpkCjwKizB
QkRMfrl/nHrRbE3eFcRiDsJ2JJEjoj6Pyh4DPHHBwwuLf+OwVBuC776ZnKWOm6iBCskfA2iJegda
Sc25ZIUcCBFivYx4zBl4ENvOcBCxQoqXkjdMjheOum0p1Z3YMVy2rgZetVt94RXM4Km+AkNYE4p8
JN4upc+cuNdfOtW3zsyU2L7ZHbXwezDhmfLDuhQUiYUwBC9Zq+D2we3MYGGg6upzRFS6Rf5jg4gZ
lPOxAK+w47XSdPkeo6pVbTfuPVvZqIZkdt81IQiMGzZlh93i9AJjTpH501LRuA5CRgkDmhIs6uDL
qRNJT03ARcZ6KTEFmfQRImwykok4I3E215BttWut2Y8X2HWwUWY67hI/K4b6EmsYhwSWS6SUqcwR
TG9PnLbz4Q4og1O3DJhwJJSJqGcf3MOkBKYwWRJ2jxedsH65SBRFI9RrfLwJOQ2tBHlrsrPFsCpB
y0qZH5gHlqmoXgjZ9v4LiAJv+PQfRVF0BOSaKFN7rdHRVoMniFnufp/KPKXMNYygEREAC9Ey+57J
uTIo5QdJgk0GnpBhlNBzwEDHnNqHDnHHBTLLctvO7XGudgW1FwUPbSCGnakVzfAznwHctWRwylpy
MekTX2tkzm4WQKbBkC9KZxDt7JLh6r0sA0J7vA/0+f1pb2e6hgQPb0+tHNCbkHaJXlSlRrBcuKVN
OPnD7fQ9ANDxPDWpu99iCBRq4c/u6OUUgfehIupHzkTgI1Naeup528wyKa7Lbia4WqJR+nNz+vfk
WV2yJeI50S8uvELn6aqcwtH9995Meu8rowAQKb5Vr0eJt2/+IHNKrf1Hyy1xnovJDndDOYBtkC/z
Z4fWdRiDXfBq8xFj4raOYq0WUAcHIGMPqlw5LmliiK/Nw8XFFUN1BJsFnmTcPOQA+7bTKrXkw5+B
sQkH/DxK4SAnAYj+BCZAuJsTI2f7+XfOdtGYDNxfqREHqABS5o5Or5A8NlZg8xuc0sC8/od4GWqR
gk4K5lfZG44On+eqMPNUIpLs3ep6Y9lK/2r6VNaGCBqHB6CO5b7ad4b6ySz7joRq4B0EEuVRXsfk
iN6JjvPPYtEA7nQ0qZfFOxB56tFBKE46qbzPgJcKt+FrB0TNbmVTV6AkL9829uov3hVC79Lnmgfm
zbdcDjxYfJEbdLa2bT9gB27VfD8cUhg3+qSwCuflZv5ipHKxyQI15ncuEdMLBz66UYPZCSAkoC0u
TLP1V/UT+P705s3oXePr7vdz0QSwlUKCRr2ZlIQVyrS+PNOj3QDMHFISsbPdwt05GGBJGBZGfgRc
0C2QxTFQxQtZoSoYjZj4WY+kbp1cTn7nEwt3xbJgq4VTbL5jW3wA2MIyvveTYJ/0pY/Mhi6KxtAe
HAp+odc1hogLdp8Vxg2U1EeocWCkaLiLi+FYT51iWplcpZdNy8rS5tuWEYDF7W1qFZ1au+A3/FJm
wnGuEvN1fbNNOoaILxGDa7PIVUbsHmNVGqA77o95yjheS03O8hDc5MFAOLULg8DHT/qm8zgOx1pK
sYYg8PwiJj1rwaiFr+OxQvviI7VP+8HP+OvMgukCuS7y3PMjQxxmlJY+7WMZzfiVGjrYilbwqvB6
1ayuKO5fASK1HD801T8Po8ZlPYixqqfBmjShCE7mBjTq4uXAF4C+4F2w3Bv1RHoMZ5lVJurSQfUH
Q6Rnm/akNyYIHMLKgD8WtDjbm788vnhXep/iKiv7BgxWXjXS0COfNB8Wo1tbZMfDLy9Wz1xhvlzK
OuDg8W4SszmGfZreUL01rzi4HpECTcDbRXhnyEy7mx6Gk7GbSg0WwyWQ8/Es7ZjTBxvlGpVI2V/M
tAcq95d5lvi2XOhTJkhUsE6B73qh7e+Z1aikum+rHxfpnGQPWUYcoRHuS6k1X2kurUoMCbdKyYTK
hWr2115/im6VsA/2t6o41Pz5DP5pxVEDDjZP23vRa31LXs+QgFLkVws32lmtekbcNxpqgsk3BvK/
NY5Cjn2C6II6eTZRHedVZ4ZkHdX8ZLvbIg82u+xjXbfikAT6rPUXtlSqLlJRf0LCCU2Vs4OjB/Nl
/ojitZMtycIRRhyzTMTNPI0nB0h3puq9CUQwTw1HPC9pzql8Epbs7Yvr/SnapkMjTLX75BqJbEUk
L2yB8C645DcnqQwRpRzai6CFprHlbuDlujPlGVbeFssTuxgfSNsiwH4aQ/OONggiSdLLJ+Cu3nSr
4OYsewrvUlPEmj/rQfegeDYX0QdkD8WxrdNKJ0Hsxq4mzer61le+E7BK1zir3+yjzal3rCvZiMzE
5CH4dgt3It5isrnJRK9lrguWb3tbSGgvUDJ1KksPLWj51sOIpuukiwtE81k0F9sAyh39wCHSGT0t
QgGOgp4mSvnQEwqu2BLCauih9kgKflLz1RaAQ3FuajLf+AiGxxHskMYEcFEUI4ZngDcVkF5w0VqA
axVJbxgAYQdEZhIXkejVEo32/NqDMmvWbRK9eSyTPdJW/Wa+CoK0QmqTT5WxDXjgvNntwgtG/uNt
fMZAfCgKbk/fYPO5ljUvlmnXW2qd6ASy710RbuWgy4WBtEUIiiW4VkUZFtBAsQGpyL5TCHjEdA6L
8LDaPZm4u2xttIZz5RO+osmiqOzdiqrCYDxPQeHjI4HsJMpz1om9z39vMhKzpMagBpB0oTF4qhIj
x+05edxMci9bLCBGOU9wS2QgB8L/m7+3JwlxMeJxjxI81X6QvJj16mV7DwDqP2eV8l0XC9j2B5JH
yU72W0PmztMznViqd/wy/lRnbF0R7rEB459t4n+RfePD4ljTG+tFHVaT9cYq7DlEjnc84NGz1U19
4KXTCIAg8JZ4W8DZW/Q47vvv9Dg4XoluDm6cu5VEUpnS9N7Oftr4izuNKlRdE3D/XFN/GDtIZMiB
MwaervpUZttjf+qoYE6MBTlPAyjIDgOHrwwluX4Au8mJ0SZBqDirKJqyOhL2BYKhohePXkeJpHTj
1w0kG4jSzQqLf1ZL55cpxrTSeKOEOMuMuALURMuLHCmZPAONsQtJBLfuGJYH87r6Qx0zZW/XCnAZ
B6VHX/By5PoxUSEQzyZiWTaO+ZjmhAvlKzEIkYzyyBVIQRlzTJLdbcBgaGhWWGJQtt1LaQaUWVVJ
sS/zWB+MCt8OOzkES0L70A7ra9i3CAar82glYhNVRv/f2K8TiCmhiY6y8VqKTUd7wtvSsSIQU7CV
6UBUwUv0dwb+o2XUWfi6/lc9U0NRzrZfRDO+O6fNFIcYg7cRP3AAVIGpeEQiiRZqMFqOgPDMBgmk
y8/U3EfEhufSfkmFOEEdG/Rbk9Vc9JbIYm2FZjA0sdvWkkMHQGcK0eLTWfWHI1h8vsk7R5cQ7NDv
1H7ndUYePRon2/o1CjHev4tPdK3SaznSKKcQpzRIrurr8EiP2fe4Xt6+HcfQLR4NhCK04/8tFDmS
/i7nt90F4oOy7GIPH9gfFVyCbjG+g40z7PXhR4pnbDmw3y2NsagumF4/H+zh5GxAIHzFu8q0RRWD
QNDaoX23YHp313EzOziLsYoatFK/9T3DWwDjYzE9JKjqhqe6uJoDhGqGuhDKIoJsKF67pASchuYr
rRTdDmb/jYYS89iGs30bKQUrHvjY3bvwf13hZcWb4ZbT7fCEIlSTsCzAClMRbYHpGsKji8mTIcco
aNhyUV356QUAmO8NnMOwAdLg2br/Xy3GpUYkZ5bue6bEW/hObkxh9AQMo4BROMErFXcMhw07OFB3
5lMBJy17NdBAr9G3NTLNP7S5D+uZTExn1W2pZbk0fO0z2OV2lsNAjilviydNpmBlFG59H5jcjZ+x
NUGfSCBIrgp2UUiR9rRoqEVMI3XSgASNxygI9f6TnCimMkK38DvztysF9dr05Z/oFBoPVDEwxr68
shK3qWEiNJWOpnyWokQIUg17gsw3UBxCoL4bLzVGRa6+36mo0H/mcu8NhrPpRV+I8PZgQH6AJjXZ
o2UdcxHHuS7ipUvAqPGzL0YzwKLFNI4naZDjHkwAKt6Xv9V4lTsnreTaAXLMT5XXw9BGU65zX+2u
bF3J36W14teV4eEPU81/UaAYQzVECDC9bJSZwBFij4BczA08mQCfYAEI38g9VrQ3NJOF9ytl1bY9
E5SNedhVTTtj5lo6Wr3JQfhuC04+MCZrtF+i+FKYXgnsY7mcJs1wr5wh2mtOyOjydUhyCtO/lj/8
gqcLAPjdd4HVwRvCnjibFOAobhcAJaaCMiqUPc57jPAF9tJs3v8xKct9HB8r6TtP9I5BNN0PV7+x
zIjx2PlVsI2FXO3sJ207CCE79EBcEDWfy3ermyKz78dHjGOMKZ+zySa7Zb2HT1tKUNpJWnGn375W
FIm41EAQVctfFiNAMbqgN5s1b4/kVsVG+NjhoOgoN2A1//zsNkajuJVlqKKxKLq1gUSUZao4rcNd
xI4Xe07Y1q+eJn951CGb5bdNc9lRftIIK4z0HSP5OGHyd4D2AdGt222R+MzjY4a/7/j4ckKEPA3u
W+ZZTdr/TAR51iCxKsE5uZiwMRtPr3ZXCIhIsfhTL61WWfQFTeF5HWdjw4Ss5fR4CYoDM3/q06zh
SmTOyc9ke4GWkS1mO0LL8Er2yQWGQE/MyRY//k6OApPFEErDv96TDdqMWZuL6CdxX7S3X3oM/hv7
4vHR0Y/dLQM/keLGHSJ66kaXVRo7E90qgV00wc/rPOtteiHUhv5O3PHm5cKe4b4Qjuas/XyRcua0
UUE/qMs26TQmgGJrfO753Fix+YhrsC3Pg31TvQWK50Wvz0uwDJt3pqCVh3SrZBZ3wajHjl3AuBRr
ypw2ku4JXBgIwais4UlDY4ZBajRz+DlBQ8Ocrvd5OuHRAofuXQss/vW53rzEVpQBqwOPnmZJtUKk
Nw6HBwZ4dY9gGtQh/261ikCzVGE1yzgjNzqnd2fxLPbYy+EVWdppIPrXa0D0KQoriy+t/yqpujDe
VfaC9LwCK4amNZohM8s0ChMgn4i22RCienhs8TCShcyxcmBg+JVyezDVZa9BJZ0YpFcu7oFeVNBJ
XGIF4TXBTOjHHxRycxQwbt+F9jIGTpjksyjzalcngeyj7yiWi2IAsAeoRLVVYN6QcaRVXSO0pPSp
CvWkw6bDcXnRtcwYe+YYDxWJI84VhgoGtMu4QqIhigntz2Qhy4ROOg7hL2KSRkk5/J7chhYGgWUL
MNm0xEP+dNh4NB5CKHyQ65LS6TeOpLypOlYuB9YNp8klWQ03fdMEnRCFq5ZWPRMNFKhu6zmSxgcV
GdOCrrTxy6+f1MKcguAea+QcyVQTsfTYj7Ton4FCB+KPRrI7TZO3wlSEqVa+HtBmCfseIzBkEEuz
83VOMJUput5sGLeokWrf3HPQPujB2l3vizCiNop6DYD+gSl4gWq9t09evGTwzUzMB+hQ6f3ekfGr
31EpVg3Rqv/V9PCQXl8MCmyNBJ4/FeqMja1pRXdPK/gerq9VT3GzTPuzOdIi/gXJCm1ML9QYKITk
K60Q8xtK5uI7vYRfgTBfH667tA7uwYBbnCohF1olHT2zPL/9gAjVyvJkzhEEyvnTvy8OpMwvT3AY
1qpYQgguyHWjhWMYGyYgd/nwS3HLzPmv8yIZe2BwMvs14R/fQsFh5qyjpYgw+rlPqtOI5PMiEpPZ
UJYF1sslQtd3HCbiDNt865cDWKHbU+iUdQRINqjUwCYR8yo7gBsUAIsSeM0aCrACYoyDMd7mO2m6
vhSDQ2Z+07lDYk+UvzOjmFe2rvxP7sl15gPEI4EadQg9bb/EDV8VFLM3qt6Ivx5bWqpx9N6L7gfk
r/X0XykHQSh4OKe1SRLjXdZyGQuj0jQZKTerMIQZePsnorYGTO0pz3rjnaTEU6ueKn9fASrky7yc
M75t58gzvuVd0HmBUyf8IYH5kxT9xdAUBNpURXLam34zTNvf2mZurSrdyroX4E/WKfq0tsu8HWQw
b3KJv/g2NpD7YExBC3UCLVsEQiMym88p5Qp6X9CrhxtaMb6h9WstZfRbXrVqmyCSh+3ixqrloCoW
NE3ylWOh6SLLwqm6sVCtsC7ruUGUFjVwRSjgbv2XKTbvIRjhLOjqC+gCUmez44vA8hyZb1v5gGMJ
a85X4cgf0PqgI0ozo4dnzHF4BZ0jiF2Gg7DbFKWQE7syJOTl3ovIeTXpnXzXIShsEwoGGmJr1cZe
gAsbIzZFYf02dQEWu/UUrWQjtxlhdZfrKBvH+qWHKA46PasvQRQUP5bhXxG6Puavoy/EZa7Vay8r
qjl2v6c6I2bfqJSSK4ey70O93vDylDRjXKdFFAsHtzM6sUYbAAol8SjPau+Mi5snLQe97+JX2HfH
Ce67YvZLsQaOVvDmtVvBaQnxKJdgjqPB2TeFpBeu+K8V37gHs0U4O2kFKq9mKLkqtKgROFQw11Yx
fq/lvcjaxmDIBBUmVt9DqYIijTSjysUdGA==
`protect end_protected
