`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Do1rO2c5wPIkTDsOW7OLHLo4j6YzfTkKqkEKT1nNoZ4SKZMwxTOA1ag4di3GqyWAxndbgQdQ03KR
xvvYfSME6w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lrS7YE05ZR4qGM490L/rpbUZV5st6Aj1ehu3Yv6Su6pEjwzAzM4Ll1KY223UxCNUJOuB1Gk8C2va
4kkhP9QeslS7hltcGZVkE8MCnif68mPbOPImaTgGNxzoof6hZ99Ktmj6wMsTqzNhFrtQ9e5bKnBo
YnFqbJ4PhKuBMw/ltxY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ca1TtQ6/884P9m3D5eRKTeE064Nd6EUU0pFpIqodrqHkHCrOvUvQHsoUPAurFiuYcqd5vkAq//zU
QadZMfMkWANIShylDLuMuF5EQBP4ojuKzBM5ePXa3di2aBW95bN5TZBLdZupEM6WMCXqL1y6P6lA
oZkmFmMQOOe5nLj5Hk8SvhaVA7DbN+qhts8S8n+hr87BFjzm8khszKAixA2623ulONYHYxuQG9rY
0I8QgXqqztuMa1AylcbY3vPn7OGr9G6YSEWXs56RAq6Ku6wNj8Phli5ylCsT/5XohdLSqMFG1Qx+
NKiV2njxdZUK2CayKQpLCPqcT3WhFuNi8xOTsg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P07S7qXU0u6S3tw55IySe1oMFh9wTBH+oHfwjy6BbJORPiiDQjMqw1cREwxtFCBA4BvBnpMCNO8r
Z2cVwCrNXVYJmHAZFnXpeyJcN503tZwshNoYmAugdoQk4JTfNw8qx//+/JGecFBrTtxK2/vaBQ40
W3T2iA95br/1E1aXp7oCt3ej4aDxL2pgJnEzO4wfLFfFW4vhIUnZT6xVa1kO8T8JsPOIyVxLyAh+
IT3xJRaNiuyYSeivKKMMrwc+Hm2SPDmuwS4iTg5tEBQxiOb29x0nYCHUd0l9D6zZ3oVZppTSFERC
3yt13kIT9DHso3JMLKChiEqPlMjLvxX41FXo4g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ij8aWT2KAsI9E4dMvJpG6GdTGv+wUF+YbVXm8oDr3aJKfSOj7DYlqMH89T6p2lIdOLVMiREWKh4J
Xo475NGlrD9PZGTE3cPgnR2IqLZKe952fC7Cc81FLBsc+CSI5RyOKbCifkY9i/8uLAnCZ4es0rdU
kUrP1029v0vCSFv4ZG3pEiEIQV1m0JKRrU3jANW54l6AIGFPZTMVtX9/6olHHzHn0oLjWWhYjoCk
3os7QWOKkcqxC9zkWtnSOgqcnIFyi1M3vSgrKhWhIXVQkfHBpMqXX68aahLwEU1hv21Ry5cYbPb7
QAxLi8ZHPi3ZkxBVg3CdxFp5gZneE2PSxOLxfQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oxyZvTqQr9uqmwIR6iNkne9JP9bmJNM6cn/MvjtyXri+EFftL9Ieyx2s2/Lzac+Homl/BRNcBBYl
1dKGt+g5osq/5XNCfmVYB8I35YM1s+kVSkw2TLaVzZ8DVkw6Zp7qTXc4szTU+Q+f1sKdvoTMa8YA
YsAOx0UfXenrgnaaWJE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yp7Mi7u4sYLm/InEfyle30/Ffcm0UkNDR7EdKiLwwxttwbJesAlS3rSOmV9BePLyOLqHLf0/DooB
baT6gVWiu5UHSF3wSFGKnjkdY7AUTGk7XPJSv9afer569FYIP6gIMc+LTm96oEUZYpobfvElC2ik
pqqVAfg07wsy49XwsSAzb3MwIXZnmcaqKCIws5vI0pmbs8OxtPyXRenyC7qhK8FYLWO1Ong0wecj
Blk9GgWZfKjkwDrpo87YOvOsTzKPdZcMNUr8t10nHDYAi3mkTUruUPnctXOZmex5jEtY8zxWWl2i
mdiXc5bF0IjD6K/wINDE3PzCMqJO5e/tNUhUyA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 134944)
`protect data_block
dY7BRYi9NGjs0QGeKUedPr35i87g3e8LCePzcLsqeXGMfPiLhCqfPGw1kiLKb3jCh3LalEqwoznC
mPn9tEdy+EF6PhoERyD71kxD+7DH0lZYOJ3gQkYg5XdcUDGuONlSRqVRjQZ1PV1zYxCcxAPzPpFn
mwdCL88QmCnfG97tZbFC7rLlWpHCVxPhrUWjmgCavtlablFbAn8k7hCDJKxmOzwW73us5aTURVby
UhJyplqJOTc7TThdwghH8Tflro6/Af6Av6xdZxkQPHd+wZ0HQCF6GlFIFECmfqp0Qf+NpMp3bO4e
cfOJLLOhfxpndtIoktYSh0iUQiaVAx/iOUUdN3e2WNbVzJEGzGmwRv7WSXgy5ZA2v2Pq2ikvgGCb
BvYl/J4d0DI7LyxrYamJ9uRz6USSzX6cUyg/zbdHykXxIphmca1uxjf3bUlbl8Fo850H9w/JiVtt
0/O4gTHtTL46QP3W/p2oK9sETQn5E0IRAA3j+449R3ABlEVvDMuK7JShCJDIr/WlYdbh9bgFATph
G0v0Efi4LoUTc0j14LfUzNPrnKgOLAOkyIbSWaTdEHZT/aoWrfRiHE3Lu1YxRDpbZxzl9EBO1S+s
BnRwiWQGzor7PAI2iVK4uIL6g/uxH6sr/aksCObUwSEs3xhMyvOvwaZFgw/cZar7SZ5vACXTJeci
S4ORpEipiNQZxlQyrvqYOSRRYIgcw5VsnK98Te4tPiqJJlTtl8ffOwgH9Iv6mld1+kyAVfj9U7o8
aBqud+PW+H/um+lAkeHQjUGbyAS0k65fbghjUBVWP4w58iO/4HzHd2UXQ6IvUhc1lbGdUZ636RDK
Kj69lWCJUs9EkZ325g21zSc6OhRozySd4iFKiMvTLrLhbJhXeRW1/BGT3L7CSGzaUMD5U/anJTn8
cs58vlOOtV/DqGo7UFpWZn9487dD/SWIjnNDTBuMWTtCKGyJU2NlE5YKgp0T9UqGflc5IOZwkLwf
71TFe5yV0roA7KWYec7+fBvoOvjO5BIGowafXh2ULETB/1EYOJ4HSqQKnoWxLH9WNObpqEtf/Sjw
NOtS05jd8tjnK1qWGuDJT/O3zC3E9m1vQJX8hZeHlUcm/9ZxHwhllXJ4ZpWZzvzJdSqJamZwCyHe
4SbR2RJ9/SQ+hlwGNVq0/WWtAAGhwloVpM3IymtQ7LSOcZulTBjox7UtmPcJ/dR/NX9BQJikiIJF
UfYeWWGS/rj9jd0G38aMsUs2mCwODqtKUXp7tn7FZlhdBoAO5XLFWlnpuj97+jKMD5iAS47NRGSz
xB2GsDCHgHLj2QFzjkD+C+iw7B2or5K8CFb84/jAUi6w0peWrbXNsQwi5TZWz6uo1rq6Jd4pA1Yj
uGk8GmU4mBNiFGHBfR7qTIx1oS52FoZD+IKgGNedKKmnSX9IczSQa7YYpz8LuMD0E5xmSlAAdpw6
st6Oi5cCLILRVYSP7B1nLn2xX5YFr8MotU+ZESFKR9MOTAxIE/oQNT8xvF4d1eHljX0YAR3yREQv
rCinIHdZSwBMC+7w2jKKImJkA7Wy/KtuqYjVPJiL0EKdXfp4qce0G5miDDDgsDXQoDlujQdKMErk
rnFNoizhr3rcy8KvKvXsAIW3F0OOMqJRFqPvpuxCOppbS3wrp0kFBI34s6xGjohAzmMVGv3gEjS8
sYwUlp5X6vUYXNrP+2KYLBCN7rKbgqCuy1NmjMzB0St/2JDs9IxD5GUERI4ah30FVllnxh2oNkVo
AVPm2ZA02YOvIfT6GcYKiB0FIsOQ3E5mcaaQSTT6PeosCwW3h8SvjClJiCrtk9+iN/tu9FeBc94A
VWKPKk2NUKGN2RlRFexA6o6zO1iiJ0S1etwu8hHkFLq+dOF++2AkyL78luhAAgLF4UrcOJIHZ3+b
sWNmX1yeppy95SlzpchThM3ewJSH074Yi5Fdwzs0RwrjGWx9ILAFwxwdn9UuoLSFcb5ML7F2Ww85
C2sswJoBeKmc/nIR7UCP7Kf1Cspg8dKKwPZjC/Hm0yoTv/EkystQlAB4tF0vHFgBRgZ2SMgNOCja
G36GqzZRprJUWDc/xsbqZOSymvPoLsJQiZ1gKHZi+qUIx1Lf/BiX71eQWDvE56/Avqzkc+RwihE0
H0UsMaxFx21FcSawExSTFIMs11v0AhXLZxcIHOERfP+Or3U45WEm7wJlBBp4A+JgocrelJG4KCWV
70YsZtELdC6uiVEFoSgmgzJB5L9c829lvlJWFp4I/1rcEersMEPP2MDsy48RbJ66Jb2EZatyHsP4
AoDpZhmnL9ucWaMKUa9raPc8lGIrK39DN6iyONkYxVCLF+IBcJGeNcJHxmz/GLsULjbBDWI59QQw
KHS3/7WXP/wstYgsFcxWDElIHlIofZAz840lV8pFQZqqz0mkIe3I4J8wO3iZwM8WWAkim8wfE0lK
+WI19qjBfWQZokAs1uPUrNMMK0mH87oL7kQ47S2xEuUnFuosIt8NvMZ5TtSHcTjND5RLFIuDFHoT
QZ+G8xQMFmmtOAcLbTyg4Jc0RdM86+7rDYZARXsmBMwtUXI+qgFLGBjQ0YmQiRB0DFshPaLTiJOr
wrlf97Jk9dtH70IEkxgTF99FOrCQgfpmO5ECMQ47r2/VxfmZ6c6177ltzv7zdCFznW0anPIK7h0+
FwOKxoiR8Li3/5cQxtNdCXrhcuZAGmfYfJRJwP9TcKj3M6daY2JbwwKbEhXlM4FF5UaYQWQBHBMp
R2mfHh8g6poIM+lkJeD2yfaLap3roQdeM+Hb9gVoNn5RURn7dy+9jukZ3FydTpNJQkMTngI41FxQ
f7ImN7V3A+i5+DJfOVdOXAh2wzRIUdQH+fbHdGPLM72uIx+5w0ZRnIh0x26qVzVKuUiJUGyn8TXF
7z2uqxLdsKOCxqjXhS3eJ7kNff0rmXN3ohiH24tnm4PcsdXKmC5NKa4QXRjcYpRMmzJ6NVyI6i0K
ROwTPyAugJUbU/EKHqRtEzKSgbl58JYzgACcKBrBCT7vtaT+bp5A/ngFcuZhEo4TdY9baWiP4BcR
y5sT9hGuIh1K2XGEu0jHdMY/3Qjc4dNzCcJacyaAkQ1rGji7kh9DMIZanJdByTZZDwNSymtonecN
ybTl66qVVoA4eP5x+rkI94STXpWQdd6iUPwHQsH9k1hLJQ4dKEHTnzoe5Z3N6eCZlZRvKcVbaCp9
6B2Dehc6TKzKW+zkcy+2vPLaWCr/fAXYdmpPMqVAW0qbIydFc+6zcaqpI+OIfaWb+ZmrTp1bqPlh
bnQs6i4Gg/FDldGuvlyFMc6/2mNwGpQOuJUUsaUDZXHPq/lNwC/3tXhdFwiPBySXZic9V7Fz7Wi/
oh5onyGqBV7KYEETyWkCxrmDAAx6dTOlav9IS/E8/DoRwaywoNNY+RToPCKZGv+ZrK6CSti+/skl
C/OCprXzzYNHY6A3WiT3Z7qqvvSU++GL26I0SL5sLaTQfKHs33rh+bxRA9UVai5SxFEv8PUeFU7O
sfRBit8hPuxudVjxgLln7kNvgoS7JfbBD/T3aH6GTJfV+Mv65y/ZkLHyLow4YTEgBt/G1+/M3ktQ
IxIiTSOtKiPbS8IhbuBuEKxeXFgXuHFqYJrnq7EC7GjbL8lbVfBgq0EP9pkVow576jTOPLDsxp+G
whVI+hSwRTVhfHBjC7MLrIYj6kSQ7aiDd4C03esHPxCgV7MFuk6fbSpwTBXVBD5WES0ByGOG94p6
uCa5fcG5ZWnKb1XFkTFlaqgDeuyHc4RWH77o89KfucqkgBO+hPNrHp1KOPrxpzimqnt3xDjCYYwb
DAXEPA/cL/LAQ6B/3nZq4VAOwShz9V+NdgDWvNl0gfmOvheIQ9MzE6ITmR9bGJTROPFbqE6JbKgv
k33NQweddDW6RPwT2yRztDkqcRJYdbBRho9iFMwsfEBY9EEEDZDd5uUcRaHYmHu4+n+hEkrWG4GF
0DStGY5oJG9wx9OEi7cLKcfXpjEC5KYB/nmcmASJpjl+42lrt8pKmyM/mbg0AJAI+SEkdkxz+m/j
M0KUn7ksXasGQfeCdLaGHa+uNeZ7q3Rjw69mYc5yQdDPEF4dYpegpb/mIN8LjVKfrjOFtuz99PcE
1lvP/BF9xmc1/lfncqDkPS5jx38Z3e5hgMB2UoVp/MZs3VKHXj5Iv9j4+I655e+IqOQSoCUve7KX
BTCBcl4gJb8NJJnqindQTwdiTTlI/IZYo5Uba1+9SJaSrdP5OjpGYhPG2nz7xpemmPsGxYxMEP/e
X9dCyvirKk6qRhxJeEVRM2iIvHctG7cM7twyvHtu8FefjLHWRGOawKfSHizphA5z9A9cbLdQvdyl
F/dpUWj7vpRHJMfk7MBUYBpSkeyme5xBqHP/DMnd+IsaH0iJaUtD1znVN//R3C8i55A6dhnVqZ7l
XfE41nVsrD4SwYZAJloSD3PIg7E/WZ8pYYXweUvQiB1l77b9V3xJ9sFzekIlreIuyUphx9b5O8xm
8stDfqUSWjFH530HlWV0iB0YIsCPxnF1/7MySy/YZv5YxnKugscP6gblgNUagdIHUd13Ka9G/2P/
ss11ihulaBKkWCXzOluaptHtk8IhfYmHDlG3WB6EZY1qmm8BaUthTo/ZU8noWPl/wEr0AbLrK7z1
cb4jF5S0STmzuNh+mcChsYLGE8uTgaBComjdWKTl2fjcoNrPoNHlMM2LCaj2+7335OJfct1TGm4G
B330Kqx5NTx2wazUJ6xXqO0WChjhBTYZ/EE+JZc7MxXy+4+fAuG0c+tGWP2/JqahZPEPTKUC10XL
xfMIYW8s+ylAonvVbQuaNWYRsuDpU8m6gN6iRlhu0y21FgCGhZ7IFitmrbynLeW+JwhnwXn5THFR
Wt+6Z7ghV1533hjAXGDYC+VLoF+8QWDr244ByuJZeAdlB5wFFsFfBH8+ktvZU+r0hEYingnIrC75
iSqyK0MF0O0isLMaH9+B4kPn3jrNJE2bD7NIBg84PVGczri+zPoeyDX0SQll6sIVMYu7EaT5Rck5
jVfSWVqDNNFMKZMQk2ZFffNHrPwmdtYGKhZo8Nu+dNBbL7yomc+pIm82DK3UpmhK4K475nSUFCfL
Hp7rV9xp4ttouCOlNH2BlH9bO3BItk0zGwRXSVho3f+PmSGt3PaIFqqRMtX4VWwU9memLPbVlggA
cs0JsqmgEbUFgvfbwji+WgClcU+sE6h6wS/kzF17oZxO9VwMiCNCaSJM78UpRXEUt5WoKi3KfJc0
MtvSXW0UcpRkcUgXqishMOYCW9SLQT+pIK25sAuW/dSgIqZVYuzvJPvFibFa4yJuMhKwpXsARI6U
Kf79juzSU31usONDypMcxD3PDx5j/fpY+BSewri57OEBS8htPqKtC/uL8Irq8qmK4fsbJum21Vh/
NtRLNq73u45GVfLQE+F4fNZLnOKCxDcOKonSTFTEtTK/q3g+qmz9wi5a1TsQxfRVIIuxrVTwqh+a
DNTL9SjntpMAZ6Nfp/usaWWXU4SK6FYUO1M3JtFHlGFKbX2IknJJPqZyzqB3KAEtk6so6aNd8Fk3
/r+fmLCYF4jNZqd2zqn2bOoKw9mi2QijCEMTaNn7FkMNZpadVlFj+LgM6RCyr9ye+PJu+bqrXNgY
m9Vzb9xBYeweLcgLMGnR91rJpxP0MdCh5CkeAq5j1pVexp/Tp0++mXYWnnmSL9HKVnZieeehKn64
eXZalu/IwEvD/6/PPW2L1AganVkwb95ehff/7RJCvbw64HknqrSNQBV+zr8iVY+DF9QK7/VnklAT
u5EQ0PX0zEv0kUYKv7amg5tqrFw0LI1wLi+BMw9UIO8SiqKQOUnFi+QF+mOk/y3XREP7yRFWOqCy
8tjiss/mCaUL73zj3gw69a3n5yQaKwGEOe8g7V+5oQVK/Bn9qyiVYBQR6C9kXC9P/ZL+hDkvr+CL
cIO7IrSOF5ARDIAZJHGdZB5ShzTW0pbH6UYLCJuWr+qTif3V49nfTmPUlJ5ZcG1Zy/I+0yK7SvfM
by+SZdxnavx9u30rA+Xl0crl0gY/5Oy/a4yjQ+Q/W37rSAFtYQzpQlrd5DiZsVoYwRng/pi+Qnny
WlmQ+Ah9wE7+3drThuMi9eJxnR0hE08gt/aZKuFmak4yEM+un5V0gBSQw8+vgypCG9k+ND+OqqTF
LuOiPLqfN+rTyaHF/TAcBkjkinm/gQinq56KMitJzG+zfMOe26Ezj2cPjKpGXODSnGwMKyeDBpHL
6LLgKKgO1WFfsJILWG4UJlhHMu8ilovbyp4NQVZc2HqczlpQ6i4JfhDMpGrxKzTC7lOj4Q1TwQJ8
4EvJCny6LLdglPb+EFl5tRSQYpqEE4Jkk4syyUGlWM2KcyxaEEEmZ5IvSrIz1FJRWpLrQSKQjPx4
BxHrtHPDY1PEZ4DTebJvB0Dsk+eoM7Kc+SEwquLLQ2OptivlpBb7d+amfL0BgLuxiaiTcaRtZBlB
RzRsmq2Yng3HDkkrDLVxcy1fDzuEq61On50FaJDcuESlmKMEnY305pxr0NopveQtc6bY9fluXyy2
00Sz+iWOYo7ma41BDpYWmZrVCxbKijW/Hvw3JaCs62Mv+dCu+5IAcLCNNb809CavDHHAvyXgyaDr
3WVqxFBEsXzcyldNhiwXi15bNcBnHH58PtzfsQDSipycSwWlzkWGweQ4poyK9CBoXZOLGLVJsFKS
zchhxS1xqKb3nBk141RnkaFbhdnMt9RGw2e+JtqcpWi9JiHsyfpsmENQvF6yciSPWY2/VCz9VxBn
Ow8/SZIdLhtdmkKXb9iVdTLHXjHg9bB/01fh7r5nIxJfIn9tGzfpgKgOu3WmGTWBA+spsTaAg57l
fiixQ+5esj7MVgxXX6585HDtKKxjYFe493A8unBEncLLnvTJOEdMK8oPzTtp6+gH3pCilgPyRHfd
V8v2WqO0vpG9U2IgxRUEvnhnItY9rxE+5Fo58TTWwoFDZq5/iXsGIVHgVaPJn8K9Ewp490tabGn9
aQUuLjciC/r+GGqnQnADA3bdRT2ycuWMCYTwgMDDA1COuHeKTegUtJXXKmEpBH0IZXOXysuLPPUt
CjmwG0+VxpOjPtHK9nJ1g5cHR78KLrZLidgSMt0UHM/JuiqbQeRdDtjInNeQfczWSM4jByhEd7vh
cR1JZhvRzZxGGKgXPD/NECkeU8akQyX/E5YILYNjsxBsXrLIooeT8k9xnDZumBJiDuQKxBmUVnLN
EZi2te06UJf28ScMqn6SU8+C140BWSwf8Ui2DZCRC4jogjZ//iRj5aEYLBx7w5ROKToJem5IIEZu
JA/brN3/++NeyQ1nt3fdRYOhHMTbzbcLSzkSySg92eEYoSIG1rK0PEnwWwIBTo6AN4ve4ltvjy27
ZpnnrRsQLzp3TpIR3nf5n2iMhTitJAc0EVaFT5AP5BrB7M3JEn8ML59MXeROt8bwr7IuRBWai6st
KpedYyppX75Zxo6p6sHocf6Wlf8+oJ2zNT6mRGejwPxVPJzNt57BF/6JeNdS7iZ4ZTr4CCfBUO5e
XCyqciOnMUK2zCkFm6zMFDBbb9MwaQXgPaK12KajQLr+c+rpgVYEp41MJ6g3kzHb0tM4EKWBrHSb
9Vq/r4TYzgmSh4NDtCtsyzvfPfkLoKRyUqjVdHv6dK5r4EfW/aImQOsMHd+d9FOmBVfWtG2CkQaE
WyFrJo+v9rv0mIZl4J92Vuy6dmbpIIpXQDShldkOtAaWTDGcln+N4AmiLjNpsWJX5Q5LnUXUEIHh
3d1gxVSeuMxCzxpIQwA6Y30jMwd7yac9iNtOUTvpBGsWW7Sy6L6WH/Y+dBjjqRPrcZ5TQI6uPmSM
m7jzeDdDJCojbXxLCK1QxfuZCpg4uuA7GafXRNywDHFso71fbvGABluoOMypJFsAF3YW9NXb588T
VCav1uHyafoUUkM21zJNwUYpkLdcNjg4tDjlNzQA+GzS/MstxQcUKzJDX3MfOzUHL0zr/iwxFCx4
DiuSTpyGqsNJDvUo4G+/kdBeZu8MAycg6xeBl9OT5YxO0Kn9+5moz26qqjPC9HPFMhlVI0//A557
Rn8xzry9saQoYhtEFrXjp0/PNSZIzg7tJtWFT1H0tcy9oNuCyyRYcljK/3F72GmZNRBd6/QWGis8
Rb6CpNVXEyFKJXzwwvSNrAWMrMIL5vSN3IsE+ihhjExaiL8M+f8xVAT+dTU/ccC8lVAxKmfYNQ2+
6AS/IrlcvSGtMkE6atYatGkpALz+t96660SsR2+KcZFANTN/br2gmPTO2RZEggbTVEM1PsK8IKHz
hJz6blZ+QowqNGj1j8c7G/THEW2AdAYj/0TnwT+R0qs1jeXtqAlXIusfEtokt8HTvhY0KvjLuUyX
OEArFmeOVFacWbwqjlaC835ai8GuddUwHwXkl7Vz46KzgeIEfv2QeYRv59QeeuciO70ngBKdrUcr
t4Itao8KpqLYT5+vPR0rmq41uKHRf2PHYLx7ogoks4kr09rOvOPKMBRUqceje7U5QigXcRIZ63vf
z87zGEHO0g3O+vfvjLnNPjmjeDnWh6MMYeQF8fzWfT2IsCECzaeaHKpsCQRclEDDHsPzqoGZrb0r
cppynqLR1Rs52P3Fi3U1arI1UCm7dllrzuspLzm9DE3F/NHtyS+GgfD3EcEbPKIOyplIe3WYCDBI
RCeiRf+6vQy3fKO1WL+3E9kgxzgsyfYU6Dxrd6ks+QUgffuUKz9dw488+yuGTlSl8G8m4Jx+FlqM
HWR1NXwzMW7TvcjpniCvhJ5ZDnLl2fa+4o5JvPuY4RwqT9eCTaqHzXM77hEJu2ltT+qHMJ1IcNft
6UcJ23AIM2clq2+u5FjrwowTO2W/MxaiibK3ErZIATLyiSA1jR40v7cn50bR2QOerYxpXN1f05k/
d/1+OKPVCRALC7ZBtpLZ6J/C/E3YO8g7vs6EzoWm2faEs71758WxgJzxZZjNV2N1bULk7vKCXDw8
GX7gcvvJQMlQ5WepSD6WBYjmvum4EmPceqG5J5yPgaP6413jjRsFu+AGiZ5l420XV+UFRTx7+LF9
yXyywdoAxm4MYB3NN6x6oDH2Rx0VgllSbMmWB3D8P4CJSgdO5OnJznq1ndKmVDWZC3inqkHGri7d
gQemvmlF77hA41o7cgLzKtaKANWvlJpObVjd97K8vkzolKFKEizPvaPRDl+73aW/gQ4E6VMGTGys
Drdadjgqd69SY/HYc/hDcdMJBrUn0nWkVwMmoQyOi9rKzAzrnnLtyjybtlA3k56z0weI76gE9QzF
oMV9GNoznjNIiI5DQS+x6h7yfVKXv17aVyvwdnCpyco7YyfPbLDqBZBVAd1LedG0Sj0sAzZ6EVhL
qx0oqExCRc5yWVtA+nGeVDKwppvOtWI9627Nt6Sfik2Cfv3y81fZAWhQQ29y65/t+8AOf2lc/IBX
REdq9i9t9SyQgAxDGfTjUAsoVxi85h7yE6Ehdu3zOD+JYIYKSwuvQ1bZRVgvkOtBrhLGilXLBE4h
nrrCVEWdZd3SdY1gr1YhUauZgaL33Yzn0qlz46JJqwF4/ogdeFHi0N8uYI1u9wx8P1ne4gSVQrjZ
GqCpoQnjL3LUcrZbM8SpdlCZUlYed80aMDiH4TnNPeIJaHvPZizWvMnH2zYuWnMBeS+h7CRlPsgq
nCdKZJxFteroZ/DDN7CF7GMKq/6gZfvtVp7RXjGiOqVG2BMrFGFICvYiPbJKfREqI1kDvWXkFz1o
uXXFDbsCuJRiQ6M7/wz1jse4R2/c+upTYxbZkx43EhKN6/X5ap4dZmjyQ6Ua/x1cxtcbedTjyrlH
l5wCIWcwlRxNtHRIQPckpT8JIkno78fI5ozhys1TsfZuTAWFKrxoWPHD3m4iJ5IEFT9mHYttV59h
2KSj7jRgHK6iivRmzUzoReo/iEGqchPGIAJmipBh720cvxpXtXITDu9jrgqoetmjIggXXBG94Jsg
fOogi1V+pW9u5z6qVM6UAscxy26hu25hl75lHULP8NigVzE4ifmaZ/zcyyxrKx0ZLCfhKUEYtSCY
tO5sXmSyzJza70yC/xev5vUtdH68Mro3er2hVHbvDUAbHb1nYgQBZ+YslvaGiAwXG1WlzWNHMNi6
qsTyDetnS7emBQ2JxKg1d1by+RyaO1q2jPDh8r3VfSCAw4T8yyk4KwnYQMKkifKq92UBAGRuiCsZ
ZKBu8N2MwdTHPjucKl3vjvMmWo6rOO1drSkxcAH4tv0jEwBCem0xEENOt3me3xCRwIYwL7I8vxmP
temkYCIFJbCgaf/O+E62FQV65he1ea9Pvmwas6gwrhzl2NkKiCZVqsOaui6nafJuswkvWthUk9ZK
Swm1rGbirMbjDyvLcErDPNn7dEiPlw0zPHG8gtzRyVtCgFz+Bjxti/RZw5yqCfVKVTlB7pcK2M0o
89UG15iB59cgonCqka3QDNSx64pCz7T5LSW9LmVq0nudqN83SRKQfkW001r7uXElmXhziPLTive3
yG4O5E3oqvk5E1G/ytj5ChSGek51dnDLgTM3gB6DBKk2YMG4Sf/5qJRc+8qzfGgBPUgeo4HwHnfO
EyjpxzdhOfwBCDMxHosSK/lQEZqOUscJSF2nZjWpDNywLMkiONdajxD4sNQ6L04Mp2iN3ouffC47
9EgYa3SuE9oj23C7rLcLeuj0S5CXPuBUWGx4VAoaEeeS7kU8hANA3enelnQUB7TTg8GTT2zPAhgx
7KSNPYnIvlETqlgHW4Q+Wgnnhq/svSSTrKarcRLqrLDgCRcQeSk7dnfDdDCBP80/03UXQ1CHo7ea
Bgq+1YZr9T5kxhHNMlMaYJyTzT6aJdWjtQPTmkJgSWUMy6v0aZ1UkvXW3+p+SaeU7+cC1E1Q4/L1
s25OpJBEVK5nqmbfXwB8Z78lS5zCjK8wjI39P3V8E7QLLE30yoSTdQOy86xbON+7nkQMk9evSEXs
pTRlxPH85a1X/wD5KRdS/FgAyubkHLKYBFs2vHv6SwpNNlpPdNXHzE1Iv25eV3fkgO2p5jgMEwL+
4CaN5iBj+hMxzQB+8QZ6GW/Wpw2Tqbg2URECvUPzOnEIaeSt7FxqNYrutmlww0eWujOVytjmaw2u
IP/Ghh/CvxEcfYo/cex7r/CCmaH/mrVqrEaodkuv4lpkXb3ZZHXA2ZtaUQQtbBYeNChmTs5ZrSez
0O6YbZWsWIDmOaJHq1hIMB4f/YSBHxB65rP/SPJxAooIPIrhf7PQ1cWfpd6VB2606nXFrVif6SVD
eBkaMhuUiovNg/I3a3uW7TM48UG0zN28lXi5O+zqUfb6cVWBguOBw+F72EzkcXkuvCdcHoae1twy
hv23bWOJqTpU2c+HNFJFADTivGQEu1gjZ2n+DwkFWFMEG20DR2e5gQKLS/BMFV6rJl8q9HSWtQhm
xpXBLeMdPK95BL3VsIubqpSQRdwN0f1WSXp4KkbuHs9gFMGMoOLBaEjgwfNajRf2k4PMY1czhQ41
H5+X/zHad7Yvor4IFviz9USjRyJ+EmKMZwBHQ5DzPELnMpBvl+UavyGX0u5CbsqysKt65ahUhyUB
ipBKcDdKIgCm5YN486GUxUVD0znNlkghGIAnUQhOIqGQ5opzeH54dWVG0fSMvzAIa/LDg9Nd37oQ
Rm2MJYfVa7lXAiAH4OxSsNDGavAq6eRmcBuhk/2cPy9AtcXddleXBgkaszYle4fwqM1aCMu9nG8U
XsZnxaiiDKOMsM2SlbyGSARXuq0WAmeK+v6CPBsx8hKK/vLgC0zYB7+Zl95nRf7Xm4tcgobhg5io
8lVG9iB5lfnr6uI03nO8EApBhNqMt8I/Bqy248hnFTHXreiKdu2eQBN4hAs2ovk3bmD0VxGGI3TE
XEueYlTJf89LXfFmCX7hrCSD027vAnX29GCPkaJebbi7VLAZjOUF5yYaiYCvjc6NWo1yff3xStfe
BUnXIMNKZ5WYgG4Kg8MUK5DBDifXcuVrX+e1rNWoBe5sakDVAGj/1a0mlmzkry+vytOKlMH/qQBF
5u22rK88YFJUfjloTw5Ob+CZw1Iz5emSjJGBmPiEVXfIufWb5HX5LqiCBaPJo9m7cCQ1PRud8lcy
GCEyMoeQ9CcwW3wLETqUKSlC27FYfPdK2smpRemApcP2w/BiJ4QTQLG5N5rYricWsymucq3DY5Q+
BOOyDwAPPlnUR6xTynEAJkYh2iOLa2kp2SvXt5S9RCJI+slOWnUX9juNWWWH5HxD9looKBFkA5Wq
1ZCv90TtW4MuVTdyZfsPvVQzyR1Pr0VafHql5zXVQxEPCoyCgtpTX1jhtHrTRkM7Ru+en7Y6xfNb
chDObnVIHEpmiNZr/NITPzKiWfa+SZkZI1JDu7eYxCxyHehymFFj1ZzJEaYVGvzgq5D+pH/i7iRx
yhfhhV6PjQwx+e7LisAQDkkhwAwyUt8DuGwpH+Nb58ICvkQr09lQ16LL1VuWz8qF7joKZfMAYGzi
0/ilskzmUqwODBh9RlpiWVxGfqrTkXWOEZomTkku1xRZp5qbF1WW2AO1KONthwpO1t6KpnhacLp0
8irPToDNefF26eGwh8C0FqtKFflruoIMA3KrnnSigYCS6UAFOCZvj5X89TCVbr6NS43ZfXrqB5k1
+bApEMjkTRIwl/ecp+jXLEv3WOJzqC/RhEfNVO80sBrjMvYwOVzf2yxDlrqhBLN2xUxow2KmByeQ
02jnyZk6q0csDKy7y2CvcxLXsemlEw2zHUU7mVtB0wPzKFoJAcS81wqc2w1gnB92e6f37reOQZrW
Xv5EJrHXqYUQ7XyZ1mpjmCAJR204LLAh2gBBZsCtKtsQJe41kpf3lppeCP6Flt4VDQ9DVeu3U4Bd
+1F9LLBerrmfk1qV9vSXGa6POqHwGO8zj2Jcf4IFO3B3qeFvVFJESawWMvi6bJE5XYlnpBS5O0lE
upKgBsu1eqC++rGDpCEtBih0Jt+H8oiOwmrwhNzG2CCORK5sp8TuxMZ+kVvgJRbBpM7Z9NTkJhc3
nM9BpZSh9/1/Rm4/lRWuzsDk/GWc9owjKd6p10K+LAGszRq7IZCpaXjPfKL+5TFdvdgAdgAW26xE
ELfWhqc5WuLpk8pTAFKTFW/DcwRPFTxQnidfP9B97bYb16YUlDsWEj2kIfv2b63PtFr+/LdhslY4
RnNHQYDauYpihsRKy/mkfrcjnVtVifqwdQ6AVEEupcuCOUEjPt3nygYb5U6uZ6TzZaEIcMIAKrzo
cfqOGhLWhMbs0CtuaJGe3FZ7s8tKwn7KdyfEjZLsPIXimjej/YK6Rgw3m6Y04aLdvgGW75hqgwjs
LeMWF2vowa8zBE7quQ0i48o4edL16446UfSjuEzUa6DLv7TsRR7GG0a1ErO14pR8z+VIEzHXEYcy
pLh4SNdrpypbTkamGFMNa/PyRVD4wlf9rQUBGHsEutLscSsUaC/vEVh29zmhUqnudsSV5FageY/g
IxmO/r4XZEvhC0U11pKkuMYujA/OOI1fsGOQbGEkGHK8aVQxpZNbktnm52+g0iqocj0ywSh2DcfS
WQtzeYzvsiuNBKx0SgkDYZIsPDih9/nKnVxyu6IEwxMPdZ/vzH3fxeHJ/0K11Wxq6DhuwNtYXke+
/VYsEO+JneI27aj8EW6qDlZKzy4NHFxCxQoZrhvnADzS5NTWTYN1HpCXazd0YqNdYWQNbuUquG2m
njv32tKLX0Jpnsi/TsNsV7rnQFqO3TviDxC+FP9u8q1obvM8KUdf7447f7o/7HRzfmeSW1RAvn1J
Qkiio0cS70S0kdZFb5lKsPm+5kOvRq0jOzD8LaBfLr2qTWyibrGBRe+4qGdDbnsN2Pmd5RbUDDS3
hXopIP/sXL7fq4XEbW7zpmh9BuQ9TIzp46SxhkOo+dnW3548jVPAAGMj+Zo/wLEqpM2j6PHicRPG
01JlhIk6OfIyKiquq0C2rXLV/cwMr9djSjdjza87Wy4s9ZGGBjPIaNqB+homXK/WmViHJ7rgYvvM
KPtlKO5io5bQ/MjcnGsG2mafml6l7/EGF+BNDVL5O29ZZUBxX5Ui5hmOJzLxbuXkfqkQDhMMkdOn
x7aMVhxbM4GzDRrFoVqqiXOE+GucmQeDdG7g4t/sgHV7l7fFtuygTIFudaet014r+Qmrsfd4Mor9
MVjsr1QgUy+1TWO00ENpmQpKXcj1lrwT+qiNL84z7oukKBp9QkWC36GDIy7TmL5lVQQ40SHekytg
1n+GqRICxvmpPiDPVRPw9PAzcwunHoPfJtxCYnH+oMd7Bb31qUeKtAJ8WtdYeBWQZCUK/BAmNsQ3
6d6iiAQ/SGddAs1nZyXhjtLxqlJGcYkm4WlvUxfnPuTWlIKaiW6IzCjlW9I4uS+G4XlpQJJgjBib
4+mFAeVAan4xLQxbXOuzyEZl5f4NY2yfG5XlRM3HU1ZeOFzl2yz10BYfjAa5ll2PlM0jTW7/odzS
bcH0UQp0od5lkqkQ+WgoByRs2o4DiGA1N8ZgV/uRdxuMPFZnmKXk8yAHHs0+IpXhzybz23ZZX0A6
jdh7wPUCiESQjoVwIsfJsp8JQlTXmRvjtVGleHCytbvLBsYeCUwhXOI6c2r0DijOPqVNZ8rYKw5I
H+W3y70ooJC/eoljaU84nDEoHA8nhp2Bupm05STRwsJucnM+1IjpfGQ/leuUNrtYrCKzf69uf1kB
ySGiaeNgtfHi1hhfO6xbhg1L8W4OInltksc9+QxX1WLPUvsOikIq4ovndniWfmfHEFufZcz8tsw9
oyypc4khPyQLo9TbRkWfZsW3MGF+ojjsDjT/MQg1pBgFXYKjO+LAwAqtnNUzG2g4zWp7X5VZEHnJ
kuzkoDqzOFd3V5A1W9IowYNk2p+wEXl0iJyuEw2N2gdpXf8lb95eI52Tt+mvsx/5hYnZSdXe0N0H
AqyjjikqhlqWYi3qMwlLxUtKRk0fttxPVJ+QiEhwgQw6mQaLqeAvLwcbLWCCOCmsZZxWWD13/Rg/
pNW4TzT99mqdbNPN5xShFxqbllM3DegNzSTGOCll7X8KWvK6YGmYURKkxoxGFHJ01c5Xq+voh+iI
A41A7/cS4//wj5yHamxlxpd2t9iJl08gSmbaolfChAGwA1QD99oUaOXujeu1EoUsz8nY7fn43GD3
ub72DMrR4mFOoUkz++bjJQ7u7eFKUW8hvZh/uuV73I2i4dRoSX349xd5qDC2VeWEUDVeWmMMPjCc
HnWePaZxQPOjX2usfumBY7aAXWN4/mtgZSjXH1VoFIdRlvUs/hngiJjfzLnpyM1P63ZvzyZ1LNFw
7CuuRcI+KLtw8n7HRsI92jTTGSdPlY7MmJyTuLIzhS9glprKTU50lPGPTTiQ9DAsXYGlI79Z9Onq
GIbnWbpLXi9Pmck29SlafSdIRpL0cr4R//ePEhAvHsi4x5F2lFppnPq9a8VxrKRo1zdMSGHp0LLI
ZNfg8Rd5RNRMqNG70HHUFnv7kZ9lC114pxIMUtu8hyZ/nm3qtR1yS/+0kFWQQNvMOOMyPDaTsAKj
dusxpQsleOubTm6O9PWMqJCCwnOZZMjbNLLdmixcA6gHO30uTV+xdo/VamQ5RjfGMy6GtIURwMxn
lP74Q447el0LtjfZspcddciFLvb1ZXQ/jjaRx8zFRx0/ZmpG3t4f4Nv2J1JL89FRxykHM6I/HW+1
e71T6OYYOiEGp8pPswLD1wIZVPawfrrEme4rEauZCHmrq5u5nsAVFl9RB31PrfK7i4sdja03AyB4
jOtVKzSdz0xhH1PSGGcG3RtDJ5Q7V1vpY2vjQrzHGRAgzzBYLgWBxB8akEcswQ2o+QxBCTI1kb54
ZL1UKORWuBA0+eIF5oXst/BxA27YZCFpKifD5nz02MR80SqwvbYYuGK/f0xLGAxseA2Q6ur0NqvZ
6NtUQ2e0OKbK86xdUpau1aprrCPDQQ5/aW7hfeWl+r0OyidnOQ7e7OhwjRchJgW/sLkDH5Lt9D/a
gDlm+j4OVGNHT+DwsrFiDlq3LUMYW/OlhpUUPx8pwQT4gvGZyCzWxSE/o5AyZJ0qVoAtpWWqu/uz
PCsleHyMITZdBMmn6AFQ0DMHitSH/nro1vaWHj2F/9crZYuMTPKg6pTAMCKgd21M0fmbN4cfvAKI
83sZLcbDoFRkype/2++VnEbus2UA4ScLL53lm9mb8sESMC0F5HZEBNJoIjlBIxfydhPMdgpvjLcc
0h+lFZrz543fWa/HvM5i9k9BfoDtdxFluy2JYWoJqVrvf3SM+i13Ve3C435g4EeFuf0bSVusGDCu
x9mynZPpGeh7HEZeO6wQ8JmSNWsiIo5EVKsYTSMbrgRcnXJpUfOIcDxjXC2fwYAEVxbSEK/XH2JA
ntPe8819WNYPaFnsHbjaB6V35Srfk8t7ruCeJ2aD+it/C1vquawhZmr18UEY66bEEbNKuLnZk5ro
nDZh7x6dk3t874HtitMea00r9COavYuH0AFFJ/vCQu0ZOK4Uhtch+bqfF0SB4bNVoDK0qCdN4VI5
dyZTaMamRchhTaFh4b1h4lZdfuTIj/eXH7zExkFQOYNyDLch4l2AgNgYNN8nTejxa7nMDYerLbSO
tGnaXDCiCYn41jOXoCoVReTjRHxAuPzh48Nt5chbg792PclvlI8DE+0Kiu0B39dF5uG9i5cdCePr
JhB4uOPNS7+OaSFnlcCHWSYjmGsAdjf0Yi/KHTJFoSjLrrpo7zpVxoSvvL7gVCN6HP9Hcufr7bm9
y44TEWT+UVO/LPTLMkKRvUkdM/JiYVGae/BEHLC4JJTtPu0K/LwLlWJ2ved5w+5v+7QUp9gI0zvd
JO6TNs+awe0cSn2xKtDh+ejdDUfVzWP7IfVVE1CUfK8A8lY2efmcgKYM9ugS3HiZRpdpPyZfRgjq
W7B1nTR+GLtolIIGtkkKvKe1xKBnKS1fUcc99k04jrZ8cotIlKm0JfolNqEyqOCSXbOVVTXs4aGM
02f4tCKNwDPgAwSQ4e58UBSVbPgiNB/DYlYqGbDx1EKKSgZEMHvPUlQ6Bs2NN4O4kNJjY6yv3n1h
9U0iIL6jGB7pgXMlVzFCzt8bKqvQDRamJJ5O9Dq3m5u1XCGBt5SMqvpSzjpHinOZ1cSm40OpdMWt
o9tY8dJsaeis5DnrQ/nEZVJ5W2c9JECSYCpNeGmTqoJnwwWDfj83JgX9xzK2/yZtCQYJm6knMdOa
pbr4K35QRjjGU4moRWtJUFv3/KrnZpEbTO13gd1VtpY221HrW9MdT9NhqUs6/Kl4Oh/d6Ct18Nxh
a4D5aORwlD7czNl/aOEtcwpsKuozRPB+1alRxVxQT4YZbIIedJKWMt7CB/awWgEAloVtYVkSevWU
ncPXA7lByjRN05pNQQUQ0eUca5QqsabXLy7UXAXxUzyIDsXqh0u3dB5APxQoj7qmr36F+QmLuC7e
nn41eKX3IBge6Ybt0uHpSOpKTY1B0kRjqmyziLwQqZka4Gdr8acGrSbIOqQvg2X9Qcjmv52dTdCR
mEGCl1q0FPNtQ5jUUP1aSeh6WTAoun7pB2DgW2AamLgojQKd0QDwhkSZblkqZru0jX9vEs/zduPU
SZOjCwOLm2qS0zV/OYB9OhokrdpUHRizGVaaXpSKol21MiDUdmtLezIc/nmUd1toq5ndm1Ak2HyJ
go4Jmk2xF7YwUwoyLAFTDuZIcCuhWAGA5gTXeSCj1QOofPRpI3+WJ7vVuZrU2/VzjsFXbKJz7UKK
uHcZtDTxqgiR5imvUmzJL3nO83pbPjj+CPAIY372WWvzxo845RmOqKZ0l+/Ui1hO47OsNIcSPVFO
6hLS8/Cg/sRS7+7PK/bYc3LkDMS6wgO5o3469k7ek97dHD9WMvufrRxA4mXJ707PTxLBMa9txhZD
aB1Rb8QErKxHVC626ZtHd5EaEM7LiLmljd+yw1I1oWfDh4Y/VHBgUDwyO6/pBmTas+IktAasLeFj
02WwQQkpzvkdxCUnw71vRuVzESgbMX7WxPTTPIyiFnuEVbDs/dhw339HnwHAzoGp6a4PdhKYiTYm
ijUJToxtQyJeMDQVt+eVSmEhuYWoklLHDs/jCvMNjvkcdqIYeDfIIwKLYZcnJ3nsWzz4XyNIvZ0G
mOTm+Kn1r+1GAPSbg5/b64BLPYxHmph3ntyJcYTwZe6AWwfgwBEPGeDJAXUuHtcxuiWrE5Woe02K
cOsV1AOz6qARC6wBgfHjUzYxf8l8ClwzUKt2SfHMWz6CuzKCNeLmpvwQR19732eYpmEY8rhxVrNh
HPsQefBfCEf1OaqGt9yIaoM3/bvUJURmMx3gA8FcWlWFNoQFPx2emwbYaRWt6c6pOLhoWc4sUtWI
22aL7WiZVxCdRn1m1tPDH4ny3i551MCawQn2MDR/GQFL5/7GJftkyS2P7nNgR35UvK3qfRvhLOm/
H0I8EDoIVJsTYVnz48DZ8kPZQx7NOv1vBHkE2A1XltTREUV8QTe2bJnuGhDONMwaSl2q4wPsaj0n
O6ciC9MSOYvHCNIBm8GdD04rve6uViprBaByPeUJMkpJ5Gumj8Bv12N8IQM1D/o3UkK9eW7rtlhx
amF9qWJgWgz6VoyIR+jKb5l+Fw4QuDriFcrv2oMVL+6sxhVL0n7W2fa2M9MjSipfKfGkdTX90xBK
XSsa6qYRkA8JYk2w/FcfDgzPA9baEeQ9V8G+lWGzuTiRhtlILkVznK7oG6ayNbETaJRu6JV5hTMd
DZzprGeiFyfOac8nQ3Weby4+8js/BdljohxOpfb9Mp/4bFH1dX5iFgbkwm509hOKYhoRSYQ2R15A
nDb6rKGHtglGGOpb8ciolZyZ5nBjHuqACPiBSQvMCn5Riz1mhfOyDMJDQHpEBIhua21JK/un/K+n
TSlZnVPHyq49kruVgTUxfgx+kbA4CCQYjOg2hOIgEmBhER7KKmxYoUYh4QSVsumWYVbcZ3deAann
/7jgETTbpm8f0CTOVtNylioGHHza5olEAlaENqAZ5Vwy6eTPgjRkcE8LSYn8bwPBULF0DAb4b2Nb
L3VincRmymS3XUUcySQpstGq2wORyTb8TNd9EEy9NZBDAjx/k+6MzVyFcWQlxlsfTtzWI0JkNZcE
r0cAr3pE65vDFyFmZKE/jZ7s7ALGXuxjGR6nnW79tWKv7nbeE0dCND4+UUF27flNuq+5zBFO5iat
c6NXc4XIcZPeuUzv2rn4kyF9FZEGyfeaJovTKAK6J/3CqIq2+BLjRcApQAAn87GA5+3cGpM7vdEq
Op5rh5gb/qAe3buoYzqgADTZ5cXPuu78Mfw8N1siz5cirBby875D3dp7jXQNYajIXn4bhJ/snM9T
WXW7Wvb602zy8iyMnAg6LJzsT5E+S6rN0nhGp1mwlHqWrRA4NTyqg+OGu4IDnTJwd6WaOxKbklzq
joBF49FihUM7ETZ14S/iMURjh/nzK+mDn4Q4TyeLQUioBi1B5UrovRFiG69gWFcQj/5pep2m62VI
BZUsJ2i2pLWwN9m72JwrDUmT2J+WSpM+qylppWHlJ1WkcBU2gVH3BI7Fy1QN6xdBEcBtjfKKp6Pf
uD97Ic7iyj/rYcZREpI1oUnSwrSlOKLeSYyy8k2/ez5w9tg+qG01PLzbn+jCp4v4v1UJssFTWN6G
EAj0KXa2LZtprrXEivfGHjnaTwtz3Hk5MSdA0292Sx66TDV+BrkjXw+IbQh+zgX5IyDAfE8RSjAL
+casnR3PZyeN9e7xStvNWhhzXUba9D4sBqB9J8anuQ45VRuPKr6pE0fxlx/07SK3nr4ZGZDJts0W
AdD6skp6/1vrwONf3c7apXwShWrFBKWeBcyXbnOUx8q9uwS6/kQMMSgYDx9ZQ9MNcrWBk/3REgbn
CwVe7NbuAgOTH2w7WsjxEUX9AkF5b0GG7RkP6iavJ3a0G6XkiPf7uDdSFab9q4BmbtyWjNRnMYRS
SP54j7enJUBbHHaAkMm3pCbCoEmbBaMLGIU20T0hsfLnQKEzQKrhYWdsvhB50NTM2nQGQ+/1Mu7m
IajD57VhKoVCPQ/WLFOy0SqF/sbGeU4x07SGZpUYWwOSJ6oPpKwfTCloVnb6LWwsgFo/PeCQ/KHO
YtiRaVAx3ZozszNir5ucalLEWr2jhw+7MQG3+ESaeUj3P389bxAB2cqTwa1T9LXFzaWIJ6c0D0Ui
YS3CSRvrlFm6Nr8qCxyM/LVhAj8mZeKZT/666wEOtj0A5LMhJZC/u8gVLOw657NBUQZygA5IaB4c
Yv07O7pHJAd4voaoJj1pLE3bpuBFrA6dQS5evw5Oi8dhD8ciaIJZH4unqxpr9xBlX0luxYJFap+5
LbsnK15Yoa8XMYIaRdYWc0MPO8/2NmV3BqRg/xAZAg9/r9CA8A2IjzkhGpfozUnPO/lzk8DSqEyd
tmzm8x41EKQVTVXMyb9OnbScTeax+9xZ1Q2dbJwrqp4FkhxUTS5xg5O17xtEFAD5SwIFs5I5KGoB
9cLsjfKc50vRW6ec1zByJZHVwA1HdB0tQlzxolKel3UotM0VRMvGrBaUns+t+b7MJ+lPTtjPBNGw
Jw3A7gbEgZ2PabnqhdXe/LN7F2Eldn6Zxtnpa31ngGbkvl3DGhxKw6t0EgPVm+sORxNvA3yzsVvX
eDSwk7BwoAn+ZZPYMWVDVgwPfpVHjzxev9lSBIUun6vCYWRrDFF2x4mVqeiMLnLco9qZW+p6neru
2lXLsIs7Jo3+sBRcvDxiqNvhi2Kc6hRdmvzpgW5rRaRRHaz3Ww/cBwfOPQK/fk0+FxO1pbzFy76o
eqPXK210G9BS4YCh7Pt8JHNF1aVW4RO83izM/ZjRGKfXgkjbTCUF2U3S5iZKBZq5aUH3UEE8keYW
8IzlxhnQWZRyBdOMvuIu2pwxBlZBJTWz5703A358e/JhSLxN4qXrLTYGJT32hf5wh4tNKoijwZEb
8jirWfUcqaSv8Duz6sjioClzHrAjpK2TfLtUm17vWBQ43vpkbftl6qFYnODzF/u316ddLEi3vNGu
W2QR7gqYAj4+D6bls7q6BksbYqxXYqHhbsEX0XEp1/Gz2RhmxNSKHDRDE0u4XwMdoOYgI/FVkRPu
87yNatrTANWNGMKveBlRo5D6VjAevl1uz2GE6BiS3KCrKCMv8NC/HwOB6Ke66nmP/5bDHkoDZ6gk
FdNQzVHgc1GKofXTivlqEXLGqshq/7Cy90tXKVgH0/oLs/NWbZruY3h3Y03mnnbvD7ISrEoUpunh
BArMP5YAvuJ5+Lw6oEav9858ZHURXXGdoPHvK9nH8IlRzFD5kvESZyKY0e5rXuE4By/ZRlG5t4Eq
ixVcG4q6p1MOypUwqo37Hs/u8Oby8n9Oyl627/ekm6Ns3Lyw7amgtWVih2MFH44rxQKdD7EDXQN9
rOxBKrHlwYBZHeq4QAshPbQb5OX7Uw6VwAZLvuyWmFQXlMofwnhmu71cu0BxpsMx56qaoKlHoKV6
zyTDlFYbkJrR5BS2iiN7nNrFN2e3mhWAYI3brpW0JAgdcep3FUq4grAAk9crk7jC9x9Sn1BYQZWg
OsykW6AaVhWOhKOwNIRYIYIcdmyxIkRJ1bUM8tmPc7FL8QKlysYRMXEQxxezpXbQWfzqXuTi/k6Q
t2PK7SaIcg9E4CAgoTU8Q+ZAwlpUGM5rwt9RIm0V/SE9ef9DhUOt9CSdr7UwU8gbheBNz190LiYn
qt5CYOn2ywmrR/dWmRklVNPgkTcx6rh0N53X+F+989f67BEE3zIZs2qxMZhGe36uPMGzIP6JJch5
wcl7+znAT+ge8+ZHqzM5iDEHohwyXmVRccFv0+SRipXvVB3+xk7YuRjeUgwt85jp3BOCkoQggThU
XzP5DqsggVl3FLKEeAAJP4OKUDCBvYzqxX/vlPZPmJR/ZUtKscW90YpZkC/Dk2iYM+bcIvEELovi
xTuZ1w/xn9nuiaBYuc6IodoDtFwFlsFh02w1EZD0qhSr7JXs7TMWc3IgMrZW5exDLKx5JBYxnEj7
JPb0/VFiCsnGCWE4XUZgWEzIuR02U8ZmEQiudxFPM3LdMXCgCq3NMxGTzx4ZLDX+7QWKuC6sIXaZ
YeV+/rfxmKDKX/86zRBB975Zxf6lqnfi1SUxpsakbRuq3t+SSagIwXuGfjjen+4u1mIxzx8HGtxH
47ZhSGITdsGC+jriQhK0UT7RvLzWr9JX41tz3RCaF7VP5mq8f9RFMm3axcXHse6l0AYKsJ+Utkzr
oZZ46KH60bt8Tj6uuflH2FAmfDrfLe3YrHyFlTydtfig5d46iw8Hvzouie1bWvamwXmKtzqesj8f
zANdOeQ7kRlCEPLUO9KHvYOlDCvAe7efzCmXJxVgsaaQLRri4glKjAdhstI+9WXGXj2AveCEBsRa
B9gN1/9m3dvm2oN+J0P48P42JM/FyXcpVse3sZtr44E/ivvuOIJp2XMub6oefgfeGEgpP51o5Eo8
WB5mSTyuHRArNJ6AhZrVahpWg5mEgrdilJ2lvf8RhSAn1yaof20dtVAzC9nAW4nGCksv/5luwJkv
r9yB/NUFXZqwShWl3yz0+jI9XoFY4HtFBQ5dB4/PoIhy1ZIORK3u/IJbliWZzvqmDBw9gzv20L42
sn19w3EV8misjye5HSMwpROvPwnfgBT9krWCVOOcIDb7vJG1vRdPCNVOsgQdwjM7p87/Ow+uD5TO
Bee4HPrg9+eAVmXErG8iMoiQFxmMMyEo4iSMu4ebjUQY0ROVvewFW+6p1zUWZDWFjxSZ0Au1n659
tskd/+GQ///uqk/ugW3PwlGlzYmphzASonRy9VVlj2BloU+F3T7MzfmgApHBgMTg37669E/JZGmS
F3CVfHisOYo0ndlHBB7XOMGr8Uk/z/w8XV21XGQ5vCgeTa1QIs5QWmwNg3ooZPFN9SHBvcCe5Fr7
2nrdGie/riNhJRHuYZGzj6N7G0TygV5Q4nvKLhGoxqjUfXnBeW4wSZ8K2LUxj9jl64p1L2TDA5Qb
lJF25hb2l1MWQxwMQrpHf8jf59f7Kj6bndanrDx6vwMnYHQ1C6pA9c3bpSpbI+ZTNVRAJA5JL1Y1
UNkz3D/9sE80pET46gCPGkb7MVWAF+hAGdw2YcqSxSEjSi2ny/I4PO0hk6GezDAO/+BlDJBVD3NA
gkJUsc8TvVbr1VTGXwiGij1DhLT+i0DKCAOJ7rTl8SGdeh3OnEgvEiiKyEwh9m2tLyQGqvV7XQTv
QEZFa1WzSB42UlCUb8Z/SMX4uaKeCqZ+rYYglbBdhZ5An6YhBFn530Ru0xc98DJeP2aOdiT+jtOq
AQKPLqhhwFRmlZjW9T2pjrg9DX9R/Tn4Wk2w0RDtZp2u94/IFsQ3HpZHXaKXo67RnbF+NALlDlIr
3mXC0M/RvNxrpkp2WMveALrgO+690sGZI6EXt67U2rSVVv7XFT9AqJxbl6JCQyvytf4wxNfSqJaI
Zy1ZLvwbvPw6UjZ3ewwFEmw/JTt+KPHMT2FarzTT4OgzTbKq8oNL4QLui7tUByDX77JKltJV/Yum
k7j4yrcTwqcyp7t+9u6JcGWETR7LR/DihQR5VdZc8475B4UPly1qnPwY4rCQOReTIkeNimYY2vV7
X/sPsZfKXQXGLYZC1XGNvvjoGL8XoELx+HunUXmdvhIIN46rm9FOjkwTqYracoK5wgbr3/+Z7Yv7
7fGwD6GvU3zNhrR5ft2uJ168fWd235/TNaokoPfg0goQhDiPagw4FEqv9vSPxzP45WlBuH29BeRt
0h2Qeo0gT1FZnXel8HNXLlAVSquWtiOxZAP0cbpjzURgXf48frqxvcjmI8H4On0qVjTGhj8P1AFb
hJJuV/UGH5XydHeU7iQG7zEfyF76gbqV9Eh+sv1ovM4AHR7kd2p0hTHqCslTbhx/H/LxMdQG1v3K
bUVusaZiol5Aapf0Sm96eHYl8JjqlfRfrgJYTwJeLI8WTWS89opcjw+ill0YvBLsvGUapsOHqHCR
0HcT/ZX1UBS0BbQ3J3zwprbeXvsi+qywoY5ymnV6qf2x5UDafacxvxarUpZINo6m8lCVuDOgU76A
XBzlwqhe8mb5nzq/+ln/kWASL4/FG3SS3O5VbfLU4Mb/qv5PpDUjCJOIQQK6v/mmeZ9tiayI+DNu
L6merECM0z7b4cMN75oIj4csEf+zswDo1SmtxGdYswq+N6Jfq/XojcNWkVh+DFM1BiR0gmBRJmsG
1Udsbi1dZHPYDPiqnV7ZNkgV978Ol2qbdETlJU8wcbDmwiqiaKnl+9XuZoCsBP2zYZTsieyjNaos
IvXULhRB8SkJltEMK9Hs02X9k9zcAZdVsoUAd/wviVTvBhqOmWnFyO9gq1jxPg5mCwZhRYiXH0KP
HAzNEx5bEGuJNM1NmjMEMAjB22OXSBB7LKqgPowkUm+JfcICm5XXEx5EWhD0M86On/S6x4Ml335q
BobIlQFsCks2xZoH8vTRcXj1W5UIOSAGI6UvDJwjQcJWI5p3sGTymEVQuru1YZZ3DGHPdx/jMg4o
NU2M4/dXkzaC7phygEf4g1+NaI6KOHAScRh6RToNxI6ckIM7Le4N5/E07vIt9JxUjj5IqZBUTxwO
YNGxXbs8jW0Rr2LR8xQMahnizsZ81EavWBOsuvw7UEMQTyl/j6q+CqI4mytMGGFPDTvnZzUNSdiY
kFubqnES4w91D9ttvu4hg7BJSdWdzfwduBaeXItWXIEo+ew/NzHTCLwMbBM9F6Biq9WVtqroZ2YY
lkkC2zUL5+PcYGnyJ6qCmeIm6mfVHVNMTdDKKxLMaq8CPsH9lqrEmNjrUghTklzq3h2D/TEwABnl
W0DIKTJDSrbg8mX5/jUjp1vNoD3ufFKusqyzM25TdHspt8Pih6htnMSFo2EHhAGpc16ZPrC5X7ld
TjQF5op3ihYgw5B6Eos8eJY/ruULw4fps5aDhWOIykus4wBjjo3j5UKeNV+UVcIOGyXiNZPdXRge
Pf7n7OWDjypQdYarDIf3r9BH/krC5fIdRfiOiqrXdFe4AZNEHOOzIYZToFkI/qEBBJSYqnKYhfWo
+VJkdTNm4BF94AAAlQg51gZmix9EbwEHCn2ORXRbKzJx4xOTA0IolaLU0/HBf6kA9A/bdlrGfJ3C
fTuh55Eet82Kn+igY38WrE66Y7THRo9AnC2NM7R0Jma0Z2Upel/v38QURIMGycNSJTQDZ/c134Gx
F4Tlc1wUmxwE7Fxnq6OXboCI+yk/yXBgL22KoJMbeQZD4c8cakdFfZSDsYL2VcbS2+bcHmO+RFNI
ysxR8b0X5ZUUUblsn1riMeJDFGgeU+tpzzriYVRpgKyGSQCHjwIa/JgCMDMfGYojI3P6AVEyUZ09
yk5P8EU+mMMkQNqoLR4D3GxOKVCKkmYwr87xGzr/zzBohiBPA/h1DSGgjm2ajKqlVzTiny3WOyhl
FEMG1atd45n6ftggToXXX69qHPs4oOBoWmqlIXAc5vk7/W9nxeXBt7W5/QzskJd3Q4tlNBUrPxqS
fGrKJEbug1CTu5wwSL1lfle588jpx1O5fxgPR4QUm+I8JVZ3TsK8Ag1q8faLVOa6yFtxP/evIGiI
ATKJvmj6lBKWAekKfj7EyCboBGjvqfi2cDY1CbYbrTUT7AbpNIJuVA84DKE9YgX2LYtA1lQbLJLU
kAa9H3ebc1GfeszSdXNxYpJ/fzSo2bCZWKd7mJA3B2UPviflkDzqv5P9n30vEsQb37mBjyc6Tucp
pVJ2xleP8tkk2hEO8M/qr/76ZuHJOJwDLfQgU39aBKq0ReTNyU2dy0dwoL1WQ8epFRaKZrjfduoY
J7VV2XAgbnsp5QrFVetLzzSDWO7g0m3bDplTfssyl9zM+cvSoP29if6w1G1iRuk4XorLXEWkjMwX
Ye9QHU6NaN5UUaibweDqOg742Lbu6LesXmz8G/aZ/vF6xgWg6FDt4aYWahnIP1vggC61pZQSBjY1
PI7GXSCxSPSo9MQOC0r+VZcuebVtYjC1Mq2kBqDarBMQeD0LJceTu/KEYcWN9VrYfwfCF8yEMQkZ
Lc+sfqqRcGMTfS0IOIFx3YXgn58JaKURjHA0hbUgzdNMxxISCew566uVxftP3x4Ny9g3J/4BBCXs
Mics6/J2/8fVm7wu56+EBK/WvQF27ksSHJwIYQ2EOeKDGMtVg7fbM9GWiYv3yWrh4raPSL0GumA2
FnMDKCGUx7eKDvZzGc7BZifE7300Ay59VGOhRBwiUYc7eZ7Q4QYLbKZ2nAUR00lakQpPKoDeTGLN
LyP8MZ49yZMbvkjXNE+pY0CbOzvELq8sW1yuEJOFB9NLeLGdRKfVpzDPutF7FTasptDkgTtSiKPE
9SnHIu7GNeuXcQNEpltZo7Pr7MSyMNOA/vfD5WnCIQr2R+uCkrpFqV9efm6YJKMiEbTvSCET92tI
AT+5yIh1pIvdrZC/C1SawOViC7L0I1gCfnHGUrSXfiBKJWUOkLFWEGKTX1XW5x3hCpsxH1GFn39u
KvYq4l1fso6ldwwrbxu1uD9iswLD43Z4FD8YMxPInInL3C2W4RyGaYTeyNmEuB6SwTkZj0Y+enIN
LIfzJ4dn8nmaf2aifo0U2wOq8hlpGmtKcTYzNWiWx1rDPpxqo5g309QEWTxejqIM+LPBeb55IVAF
ou8nbGqT7L5uqA33gQYpB42VAmyT2ZWJq3GvcBzBCBEP7B8Q/jMxLa1jVjeYWTfjyd1gDaFBetdr
zqMi1B69NvUBbMGZBoO2E7kEj/ZGsFHcibr7rYfcQrOF8/Tyf+LTjtgN/bLcmjK/oC2Vk2ChcC/0
3irCA7NBodgFhVvDj5DQmW9ftrhm24S7OvMu3CW6ViZTC7LOyuiRzBC8NE7wuLmrGRMg1YHBs3D6
ZeP7Zg5Cpyn2VWIxK9B1tvKRCDmvPZcqY3FSwWdIQkVF8SPtnFTBCwr8lXxV5i0Lxe36Z1Hx7O/8
ZOuk0rSuj5lzHyGls77jUTxphsX3r/qnSCAz1Io/IvpX6jTi4n4XGteST5Oy342cEWd+rLabcFWc
i8NfomaqsbdZmRfubrknlXeUvu1ufKSig8DdM8puhlRiQxp4Z2FF1BfyBgXywsEw3fjVc5B+iN48
6C7ujE2R1N8R0eb0FtEl+5+NG44P/bwOFdxNlOiLkGPJU9iNzRcnb3Id/JWqdrdkmwj1UQvQg0g0
nPnhJZ4qFQ/5IWvW324fdMBhqec/yG/wDwe+ii8mEBWA8sF20m01bkSHn3liHujSa63LlYCpFp5q
x6A59C7FAi3lUhG1cBMIeqCiB8bKxKDVTHQLJhOYQRju/kicKS0T9goKt+EXJu1vC09HxV8Q6acg
AlDs9Pp70sYkiRq1TN3a5S9meEeh3fi5b7Ykm+Jl861W2x1TWoKY4Ow+AIuYZoQmOY0+qpXPRAIJ
HwBIn23zEL1FL/0l8oc4fjRZAz9ZwEnCkHBBEH8ymIigtc16xsK3Akb9YHd4K8OC9LrwMoT02JEo
Jj4p4OFYG+VldflUwFaPHOTvdGzHCFgttHVW7h9rWWuDaEhdlzMhtGchtKtUtoCB6wTL6tlx0n+i
O9T5BeI8DYwv5FIzhcjH5JxHEq2O9o61IP3QJcGUicCd4qv3q+RWEeh8ndxHXPSzUMvVYJYMzB6a
AgTFsuiUY4/2kWnw6tCvtolXBkJCDx9xwUJB+tBo3tdcDWIDR6EqobpFgYbGp+xk2SsreFfyH9gh
PrWHlHrUgf+56FAOfCUxHdNYoJRlg3oShiN3LnkjQvqfQNb72k/7GGnekgK+NNDznxgGqi/psCu+
SCHAaSZOMjZlT+jCorSLa8VnEOeO1o8l4fI2Hx6zAwbHDxKhmx5yHGOxskD+3dc1FfhsH5KWovmW
GHgHUto77TX1QavBhND7jTPtTdx5InHHjTi1PWcapaxKda8qTQ0XNXCqPY1Hc51VimGPfiASp9HI
dhYGHiAAG6qRHCEMGD1N1KddwhHXGtQ1AZJFY1tkJ2QKA9Hv1OFAFwrCeOLFaDbMTIGlmWJKeMER
QrsAyE2EiR6m0RfGyIhRX6LrvjbqBavQNA991RQV0xKPiBt40Awq1NiOZm81s36cmzOMXN9Wq5uC
+2jFt9I2s9hA+OYhTQVpV2wW9KcvPcfQUzOvEWL02YItLvmTcl1NLOOYWiB0cw7A6Y1S9QYiwXiT
57XEsfQpykPGb8FY8kKlsgxaGByaw79oyoKAaTJkkkXcrj16FSYnW8D0U09lp/p3F2DuAb4kuucd
sNwFy02m5fmT/fIb5OzFDXJTbrPjxWl6tW0r5yJ5GyNZcJ15e73EHNX3a0MN1QXWA378Uh2ZnaLW
Mm0FmJJwHRJAthscB/mp9c2RQxyRZkKRfDcVs9yuoIY6KuPzNZ/VxyiVjy2oURN2NAmz10GqUUFG
BumnlRjhUvGi3Fq5meL0/FWtOdU/wBwF+tEu9cjZI6rvbUbJTqWpZf8jD9NFN3XLIM1gTiGzFOnh
ScSpi0f0ib9hladmG4I8sV7vyZlUwCGlJePeWA1SKxd2oaHtSoiKOBqGLXALMdR6Dc2sgu08IUjx
lHaZGdFT1TbbXfvyf2i+8qqRC/LAdBVoTV3N9fhUDbbopbuQTyS9chosy0NC45xUaB94oc/mg0Ae
F7HaoUiXoeeHDbq8R9ifBNUxN2wcrpo1q2qk4oJnQ6wNgwGTR3LW/eNDH6op9MWG8EpfMP/FgIHj
aZKrd44RBjpsN32g7I44/EZNLiQFddm97waYyFfxk4Sj5S6Z9qxBJP03fWGeCITdWNzFCsoGr9Rj
p216svgwMaVHtFKvf/ujjsTxgP35txYkNbmki6tS3eBVxlsMICfpFtkp86zZDriHHpAKomjNz4Tx
Cc8ndar95BkwtsqXglcBN+Kr2TgDRK9OXf9XIjCP4a6/nyFC1wri3UMf2zP1DsgJQo/N0OhNS73V
1KrLOXPKDvugG0jGYh+aHlVLo6db7c3pm3oo9YRpFDvnloWj5j73RoYqr5vfv1IN9uRJwuZ7I2Ao
TS6KHhGaq6RQIFc5q0mXwHiWzmoZ8Yq8kOsVBpuM3Ed9FzFW35QZGp3cDRCAyIEzTmaDHNPVnmvX
upR1vCLQddbeAB8jbDq7y2rf9WE/6sJkAzRAw1fGNb62BEHcVHguXY+6VFBJAcO48hinedewvvTS
/KvDi78kLAxNu7ztPDBl+h8Szrf4F5MuUNhLQjuF17qQjM7g1Pa8b5mRS9kEPnbSt9UR+eJakkzJ
112fqbkQOdZXq5WB6KzulmItcSzCyfnrlYl/05CIPtp8TO6X49Sp9T0WeymrixXjNTcb9unv9DD4
/LqojmLibbO97bC0aX1rUbchZ5Z3pjEfP0TgUkBOMLZE4pzVtG72rx9wjfuEPaFGqxckZ0Tv+qv7
9BqK9VgwJOWboOBSFjXm5qZaP3XBYPAbK5AAmLWzax6FADAhbWmZjg5I+/duhog70vQD9z12f6i2
Sdg6DuM2zwE1OWZRzKRbCf2EHd61gIdbVLdNFu7Ote6oT0ZqqSfylG6VtWKTUrKfp0h8OUBTZbJ2
DsRXqZ/HU8Rp/8ah5KvotxCrb6nYr/xnerzAqkWXTvfwmre2CArK4tAOmFofJgtM8QS7q4Kv3rGu
f/HzAU35ct3f6ZxEiXKJbr7Hf2bJ3VgxCEuG752Yh29zixekq1o5OcENjfg4n1+n2dmwaH0I4Lzj
sotuA0Wa0/nhIldleJ8zqaLAES0+j60r2JA/O1fqkcy2KN30PiejMSyZ0sfLgAuDXGzobuRqrAzc
KRvAQF7oM2PeGCjRcsGLq0pIVZ9hMTX2ktfxJ/fuXXS92918qiWHefmLAUaZG8iexXI5YPw+m77G
FI58zwmuJONeuwQiQKg58SAgLIGGOuqr0U8cheFgjzcw261kfSCFNlLBCNkgW+k2wwb7R62pSyv2
49R1VNK0lPzg4Y9ycnXclGdloantoldebbgm7/BPL8BpPsDah0sWcQYxrfoERW5p5+XMUt9tK9CF
4gmt3SFr2AjFLtza295OIjBV/JGSECmjSy5DZTVk2DAC/QNhl+5LHrv4A+vn2xf4wx+Kv43II2WO
0ayq24/A+2EHvseUg9Fkdudww35j0d5i4OmH6gtMgyiK3A7r/n/V3BHeBMNyv5RDF8dHy/Gg4J6o
EJI6Irrg4rhrC1NPaM1iqAUefwncUI6lFhA9X6kxusPgPR7ggSYrB/hPYf548HmrXI7keJ++UoeI
3tngfBXkszLV1yLeGIYB+AGz/rnTK3vfvhUadAxxnhwL/vDgiKaEVWKXuI1NW9ImyXZf5/1r656f
bVBquyNo4P3bcZ6TAUWcznik+OltQhQjTDtgDHiVGgpUSO6+87sw9RNUbcT5wSie42m2QyWjiN7L
8DY0XftymaD0K766PMlRD5uW9dUpEDlZWQ+3Ya2OeUp4O5DPW27QC5VTgZE4/LJ5Ve23DoY9QLz2
cS8McSwpoQ6QJomSGa6iUGuVt9m7SGUei7ZRaPX3p9EknuY+u0tcQQ44nvOZRcUl4Fh8DqFxSn0r
V/1Y3lDZf89Gic5piV7F6EdMEeOjDCfMNxu5jN0CeSOECFOFZWdyNdPNOwIktPVcBIoiVcrAaoV/
lbukIHwdx/0TywftPTbhi8ZrJ2YPnsO9TQgyNw1dPimv4tbiBBT0H64iguRWvtgxqW1fIUF86OdQ
yRTGPPiG9bo2FVph0KrbHzoJAB/Hr2UDWETvNie5ULtMpi/koR+uA1IBpcV7BtUDRsg1iaC86eRF
xRpkwXgaO3BDRdxTUBqd9I8tgDZOiwOtVPBI9Ow4K00shpAD7m0YYWTw/NhzkIRWb8rp7Ic5YDVY
ZhqPaOy/zz3WZPbrvhVT3l/B4+y014zsmcfvLzmdD+5rGhkTWWMDhz35kuc7uv1Q0T2t6rh27qXM
+sr88lVw7wMUfRiNSK4LqRfZFPoQU+88uUu5xEhBSWrn6qkNZmhOfIH5GkqpY4/CO9U/8mtoNBeB
P4+F+pSvg0LGfPNC9o06WeiRDbIFnIAIOlQUy/ECDhKPxFawwBUSesOVIVbvOtNj9CiJJ6GhSBl8
fSO5OP+tz4CtIxDlikHcN8bCxZFfioEfL70LcbWI4/tb/YCtl78IEQT5Bs1XbSblsBfTw78om65/
foszSMWFD+z0IfunMWemgRHLS90K0hY5ejpHUxa9MA9VSy3aUDKN0G/k7kMd7rhiKO/MZtNoNyWc
6c7pJro6ekZK4OsEir74X1BKk5Dai61o8HULwntoa9HDvJtID9LDkLtUjI8GwZLxjdLpeVQ3tAs5
18b0r2gUnkeDZvSBjvRpxwP7vWmTCQGFQVHBR4tnEKgIT/2/2uGvXADpN+OrOE2JN+A7Q9uy+Ysk
DQcVrgm+Tts+otePfKuiv8G3LU7st2HrnIajvyUT19SxmUJU52R/sL7dOX/3BjRONHUJYil54vs7
XUukWGnGVOfxROM+CT5fF7GpfiBBEOLmj1vZPfVXOFMKVJjODriN0WcI5KVclESi6r/GKjk929ex
Ts1GWeleUJ7euUi61Knu3mfTdByo0BFpJrV2JuTWURzWbd+c3LUpKAG29vl58KDNfqKTwSweCOsb
H0vsVDSK0slxwdyERM5ytGBXBCjAdkg8o+gPEEiu0yc2n4Vfea3GO18aI7W/DZFCJC0VkOjUhCpk
+IdoX8NusSlJedeTiHeEHdjUxL70XeakFgrafJ2uVrEdjFt4h747pK4DtimSW3lquUCJyP7b2CMX
YzqkWiend/UUdic7xkjjwMpzxCSMsQGHMd9//CwV14oBwfskWM4JQwVDPy3/t1RoOuDDsZGfd0ID
TveE3ctbDQkp1bw23bCys34QSafmMCVccGs9enRtQT8m7950Mz7o8WAYonRQtQHGw+LwmwcQhniT
DgzI8MsWbpHO1MwK01Hwb0bvjrxq4ZIy9IBVuPf1IK5FneoG94eESkPNhxjv1kGXOUNQGMsKDNwm
t+Mm72NlDrLhkfUp+CN/xl/5U7iPLNKi7cHPtqJXRmQSBynSalnWNh7IHWsdixTFFf5RNglHuZQK
IiL7+GR+p/NI/cbeElYBDrj90IPA1qOH4dj9TjPc5hyxeuXyHruOUpHSyt7YPPn9t5Dd7nguW2od
qDozw4bzOIN3vDMRUL7AHO488wWFpvFVCPV6HmMmY057e/cUzQCTakWaGnRbietXG1hHgErH8Mvq
rZEzzpoaMwJ1Ump+eCanOjyJMNobrayjWrqTdpM/Ejwm73ADszoPKpJTlWkRcltbx8iEETUbgtA8
/RtCP/MMUk+3FV2mrfrhPz0LuD4OVI9qwDP5hV/NR52Zrn50diTr6hD8r9T3upAdtWeU7jo3uWKR
I4xisG4ZSOl9O3PzAOq8SSZXL6NJSJGczwU9QjakiKTn9YdJv97Op5yDG8zMVDVlB5cSU+VsHpOs
7hfekvt3qgVurr6cP1P4pYFC3w5B07W1FInJsAatRD1SKGcc/JD9v6uifmIm5oGLf9fKdQT9kPcU
akJZUGvFWsSHxPQSECax3Y/fq4gPLSXmwGjzzJJ+sVsfNdQEOL9EIenVDUKlSPXK35ZqwWFmiBER
dVFsAA1vAYSfxUOPpem440z9LmBiFJv+3U42kyfycUoC5nTDf95//xYdlZrQP2kbaYoCDeY/gh/N
L8/0VVsiE4YgL20h/1rd3RiGZw/hDirJJDpIdCJyiS+oTRUG/4M1eE3VPH5O1X6qXQK8fH+ncJCB
9dOob5DsQNIrXFvWFMOZBC893vUF6GxR7EzYLui+QuiZjp9jgkkh9bGr4QtHQmvi2BjmxXoBG+fy
UJe6HC7sWEpqTx3gh4Me2vvOM8Kzexq1+hhackYQFMBvTIXf3Ruq99zIQxlSHf4OoZSp69w0wbF4
MRJ+fLhk9MmMk60FP+S+ThECMkXV1ncGGk1XOhwECm1t5uwAVTbrPL2omFaN2u+kVZMvBS/sn328
z6OwE5FLCTiS7yJizI6+WPX+mAwi1eclfOJE2QscSJQJUHgcuztNQFahNd8ZO5L6qSRl9VYTkPvi
oTPLuQUP4BgsVKLk0+FjN46DZYm2KaMCwqig9rNxeAlv6uNRRV53ljfUuRXrPrAsm9Mmu4PkYhlC
g7ID2mUIjQl71kNiHiQDzquUvPx6kXbpYAcZ4Bu17NH5k+ZFvXTaJtQUBNYek0ZIFJAeELUPHAdr
76aSEgG/pKXupCob4aeKB9+0wfQloEgnDNQU646RBTrxH46SgOxc/Q5s3VQlu10cZPGTsrZuj137
zEJzuq0u+R3UWzSB+xBIkoUJSME4gEapHjCwTscRGAseuV4AHxqCcM+4ttewIm/re6yNIZE6p+f/
d+7wNrr1ot5Kp5U+6Ii+jeXGuy19QYAcO4Ko7Uoky2u0I5a6ldxJlqMMvOtcADT2bvL3OxgAnVhl
29Kl3ZOeoY1xJcdu+849d6W8T35qmrssNa+41AZ2dAXxHlHtP4jSVsXR0z5LAfmMEBkZTPKBE7+S
VhLVhv+xntYetpaLXwoz8Znrgjccn5ZPr2xl3W2BuvX5p/abQqrL+DpqJs1Tc7OOBPHXEueCEW7j
7MJF4EFX7pYxFZL/6qBIvZOav9kZOvHxy0gyNMwajE/uq4YKagIMBRAnz7xgJenwe4caV0TIiMo3
xmG+CUKwBKfPmE0/xiztipC9KMUPYc7B23F54EvgbNrGY3/R+o3oNmQTwzMbFZpweO0+SlI6U8ez
8YJnO8iFHXjyy4DcA9QhJvjRqteshhQFUQkUTNnIUy8CFsZBGpcK4nKrZptfV9bAZ8D1o8oaR8cE
F4MNm5e138MqpJp2B9+qiOXMlChGlJVuZx1x6RfJeb5wagkCMl/AvbK+KZpshZaif1b9zHQ9+ENC
drtso47KXc9jnBzWG/lmDR58IiezNyVnE0V2nwqKFL3cfIG0EGhAo+ZunokiSebFqJwWWzIHa7N+
IxkNw3aOyVoQWg0BblpCNTry1ZAsCHUyJrqcCKy16ubaH8Cfvjgz+IxV7LUpmQ0sQmthJGPmnaLx
d9nEnxx9eEeGTJVHTGvsMFUDmoTFn+2EMD2apV6sgZM35gAfSWqV97Mchb/Xj/M+rVUJvhFBHWUA
IJxS83ne+0mdi0wqXh0bv4GCK6qc6RGYLVvEUUIKsFoFxyfRwApwJFjy64UYKrQGBVNec2Hh9G33
h7qp91caIS4w4oaWL0MqeFEGX5Br3FDCzYvRJUxTdzSQHoIS03iEYLSbihBtWFpjy5R+eqlItl/3
OUpXHVncxb0OmEtqZytq4RN5eOvM6LQMovHniXrTF75mmnHnIiwHE67zPmFl558zAzQ48E8783Fc
m4VFEvnu5Manv8ipuArTnVfW4VLiZoM58f9QYqUgqsIChwCfPAk6oVpu4hHjq9HIOOX5Mu+2xJuK
FCZjbyYh9e4eaPx6rdmDI3BGzhZxhc9g+/vJiI7gDkUx5g2qHZNgF8UBKf976oCFAXZ8qoH1vXD9
pRKsjAdZragp8XynLX/li+Grw+fvvWgauVjTf/dluCPzy9LYnmOOH0a6OsxCsC8C7JZoRs2eHKAU
FsN0L+K9AdOjpVuJqiNZhxBAqedI8yLnNZ1Owc4TGbygjIP9pUl+gzmisvx0DndsCRmeUEgFx4S6
WUAUSKtHbMuLrFp2lVxre203ggVNu4bHhKZNqoVFWfm8v9a7o7To6owsXsLoPlseo0/jeskwTwSW
IsSOxpY8kdaucGsa2ushU4vVzaYY7H5+U8iUKA0ha/mP+NADyPE66Ko3HUySE7wg3pmn8qIgbcbS
xDNISeDxxt1YXWWZCcSLFhhCUErRby4iKLBQh2iEgYobbZLcVFDzYoGeLWhbDT/TqzlmeHnlBVa5
QlIe4MLAKqBmlVYmq6qb/kKVfkl0J8oEVmnPj1Lwvd2pB2ItOZFJIxj007D4EbwUJ8fYtn54WHp4
TKY9QUHYu2IOGBvg301iQSsOZsxmE7OC11er25/6Db6jxCIlvKr7H4EMyEZZzSnyXNsKUo2B08+y
eiI1IIOXZTIYSJHukj3DDH+r0g7klb2sPUBIl6MkbxLS4ysPoJpXcpFcYWJawXJJNB9dOQQ9zvpC
zHLj6KLsEpUok1fQ+PfBRXkizse5SwCg/ag6rlrxaYxumylZqyg4hxprOGMXBr1jfxwHfJ/Jgr5m
cO4zEERlB5xwr/b7mqz3nGplL/jqnoZ3MWbOTHS2EfzxJSjEd1tT8hcdQtd/2t1ft+z94hcKpwLo
7A3MwoOrkAsqEGUvJMg1Oxk08oeeE3C6NOkUGOJU/UKMzeWd1AIbcQDksVE6D6PhdKhzQKemRa8N
pKEtVXuXY4xHPH2c2Ek8r0kZFHoFb/hVqcXp2V4p3Lx0IBunACzrXnQrCSmdpCFACLjzM62fdcfc
heE3dGzBi1JzeSbkKlRT5Iz3GEJSa+xVa3aLhXYNV0m/+7PHgs3ypaH3I96/CiYFOMW+9HOVpcMm
ec7PLlzMyXsE074LAH7qNbX2vDhqhWpwdL5nDrqqfZp56ETqccKX+JoZ8t2qxQzvG+junftg2Y1q
6PgZ0vcUgHMV0ZZcsU4p0r9ux0rFDgs0zthcpDmCTqaf9cwjUEoVVpNDcJc//DYqtycbiOreqL98
lwhFLEm9HdyUeQGgbwrUl2q5XXDk9gBPCifXzvpBwJfa/vY0G22pTWYCG9OSviiGILqeIY3GUWyL
3oceG7ShIj/OgloOTZFOaDtLafHUaSdXLX4omixL1FcSeBS7AS08v0p4Rda86v15c5+JE2rB4uSD
Uhequ5K8ARwt1ejpZsX4CNPTSgj8NDJDTws8eFMkYBbPb6/wXtEbq0RZ8cK/3EVB+PWQHJudOqaQ
KtHsk1AIQJ1K2Yk6U03geYAnRiYaYz+LSdnlVZqwkkcLEjwC7o5oESKJWlpK+Ly6pBt/gZM2gsLd
vXTIiQ3N4S/k1zfmBMvA57XPVt6jtH01S2Kid5m2WQl0BhJv15PBeUIRDlPFNGPcl00iz6g2B6Hz
emcz5WOtDMHZaW/8KmGGMZ3H9C042hL2RpmSLxxNgmzI3X0Z0ft4gaYx8gTyWABzqCpqMr535YDh
cHZ2DPAMR1xyOEJ8DXDkPXFl0N9zA7d7QTQmE5LZwUAgn0DKxoS3+KAkWZ156pt8JxZunl4ayxnz
/2Er4Vs0l7yCuhPFxpNZY7VOm+WYohhYl+rCLkYu7bIfmtwu0R5ZHnoNVTnGDZ1c+cVg0nVV/VG8
y7wZJ5er2Exrw/KAEeZPW7aifTMfahOyxrf+YJ7xMdpOWPBMmsZ+KWrQ1PsvE6B2V2nyT0ar99iU
26V68pWP4KjHE3AJYtxAo+Y9lx1vFRdtlwShQjLaQ4mDJ5BFypO0qjTbND1oUTnx9xhVby+4DCDs
naW/az+7QuKmGe+yL6BRseMy7OHd2EWP1+72kAnPM7OU0th4T26QMvsu9NeiD7O0iXanOdH/hP33
meZazftpY/iSGShemLvU+zBN+4+faksBgCLl6hDdTX9z25x44ibdL2U7boaaQiYjPU2McwILt1fw
k4Bkuh0odC52AikZYG+NjmJ5PqvBA+TPsD4icRuKXNTrU6U074BEd9KhUJdKhp0SsxWFwAbJ180A
wNa7FqpPZApIrfIP8tJF+MSgDPEbOAHxJuNDBJsLi3XiVFE07jpp1cp8Czl28rFwblUYkww28ogl
tzoZlelb52XtkeYiubmFSu9shHV+YkUCqsBCixz+oHEDBiWo/PwlWyOj+3qeAEH8RDS78+xc4zgz
LjzRmSuuZ75RxNcyt1K/sea907skQtrUJXf18zk0ghYghKT/osVbbal0aXUCyyeSpU82G/E6ycTo
onRFO07QRQKGONuv5Z9yQ9Mv6AjGYxQSD5wlhIFMrjy1NRAKnV8eUfRbBjNHK7oPO6q4Jv3JA16c
/dZxGjiAE5895bjQlsW0hDJ9KYLARUxG+4JfGx4bkjT71Snvv2UNfZ6A3S7lYjR8uMTL/jzgLJcC
8CK8vnEFMizAI1mEHQzB5yZ+XCkVbsir68TVvJjhP5Blsp7UM43MOdkYUqDoJDDv3UT3O1lzT10W
U+D0s8ya6fdvypP8Npc7r72YtLenVXNXdtWJN7ghgq8f5+0Hd/PO+7yOlMicFNaSgN5xhaf5SWDs
N+VH3Q47G8h7Mu9GxnfJ+0EURtgGzNa6rRfJJaHzJeYs0RvLRMv7H/uWLcUlaw8zAl9xjqAUiXGB
4gcc7ZA0SiZ8VFVuoKIAztXHAC1f+zBD7ui4Ia2d+e4+2gHW/wztu88yxieiYoNGjnv3yu4uWQoF
LWsSjgdsXLh8QYHNo1FbTzPp+mvM4sQmSkFYRa0BDT9quPzaijFIEm8y2CksD6wU4C/mHzsIdUW1
/aBUxlDW35slZPy4+TGDZqEUgbArvulXKZybP4mMQiHZQ+Ba2Fo+Cbbh2pid/3IOuOPCF07+pz7o
PIh+Xk3/v+IV5M0DA7JYEN1CrrweT9p1u2yFH4UzAtlkIHD/2akXZvZ8pckGW6qr9OT+753SwJUi
HGQZn62XNPcrVf2xwFoe2ZoRFBlRlL1BhQ/nJ5vxZvszBvZIvEMWgpNH3ez8g6UvVoD95aEV5zeT
QlqalgUEOYO4dFKXU7Sih8Xyl7IuqyksDQRXViT6xO0zc0Z51axEU/WCkFpAYcyAmsmxR8t+AEj0
TsHIwOnJ8VhpNwxryR8b2gu+GIzWz3Sl1gP9k1P0UYYbaJ6Z+PlbCTUztoDKdco0FXa1v434Oblr
E8nTIa6Px4LdV0f/9rLzh5vX35V3nHbTzylGjVUVbPe5RZLuUOJM1AaesyLFs5kAmLI/Z+5pJQt9
llC6hHb7nqJwUa3Vdcr/h03rDc3YOYekgDGumHv8EdsP7LUkaB7KRmx3yvbjrxp+mqtjziz+Tn0x
KLzwrlXGCh/FkwJ0w/QCcoUx5Xpsn3HtwmEZQHOYyxhUHAi+brmBYORCA00kEfi6UGKIkDT8W0Dq
CHFsh7H98eIVZQR3YjpPZOlC8y+Ec9qMGGLcxzgghZD/+JzsH6C9/KcX/0T4ABAF96kM231IIyQU
TDnrfh/QZjFMH7ilSy0CwwzyYRQCT3ckfWpjf5HEvuwdbUL0OfSIwzE+LmdJTrVm/omjDyDAYRW1
0Hk5Z0ULGzxXnggu8eqOt3Ds6u8KtsZyiUXQX2CmQbO8/M9Nn48mY6Ay8gDXYvessy9hlKEONJWs
ROXswV56zjJEBc3HrUN9vbRBEfkzBK2b93C9hBsBBl5PdbeRv63B2Y41/gksT8vmC454SX3gr4Oc
OBLDRxHFT0EfFTRivf2c/EAgDNpFSo3t8hxe8DW77jwcmThbdZ9s8ohhDcPAdaPH4FlGd/EvbIBR
GMgFfVcbR6KgqVTR653LVwFBxqzKfM1A6w/fpghO57VFxD0IqXgVLJjWTo6UFZ1G+rdFaX8OHTtJ
iFTSGV594j6Hp7r/6LmteW1bx6R21DdMG89d18RRtR1xQrUMNGfwUhynr1iy5pjSTs2ww0eVnNtx
M1dICUAbRe5/p9qB24HhXQwDzZX/OMif101MQmcEXlq6QQuucRyecSDATRDVDc3cvo3ilmzGql5a
6mUzc9OW3bD6MxiIqiWABRX7sTWGNny3+9Y3Drd+ZxlnWryCBqpIWvdlICat4cVwDxFfhBnPJM8h
LQOA8ntfdDqnbgmGIQT4k/l58B/aj9zQvTIXTIk9uej8r7e2ZKFb6Rw0BAJMw++o5peYDQnRny4B
HN2uJwRn3XtYzdx7JI6sj9HBgUe6z2chHZiSXe4oLoZnFIQjN9/XoDIefWiUX+KHQiRJbq3JqqJu
itpSGYYKRuh9bDia0LiTl01g5oEJRnnhHyKDEEaB/tcXGxCNkCEQjZPM5FOsZ71stikQIJBkfnv4
NMZwe1/8+JYC9OxC2FZpS7EFZTdO/WjBF2yFq/ovxnyR7iF8iDYLDN0kqInz4PrwjRv7wcCOSxAP
OUP8RXPgQf+hLyqZlqSC1LgJdirslQT9i5wKWF3gH3d8s8MKFP7OPZrsK372O8BKV5bEcCeXthoW
NyCMY3yY8siNZrjBVGIBfjjjEoTlNIba8StUKRHi+g8rTARfVuSh2QGIwV01sQqwS3+m58SQgCNt
oUMF5ofL4Lb7WuyZGC3FAv02idhL4LIVC6/M7JsJ6RvhukTchjySkzuyLnUXEcCx3Tg1Uj4FUH56
ZJYCdqqX3l2xi+dTgJDx5oWsc9IqQ+rGvpAphemZHmTYKq3kbwXPedPkooyIC/1gqwQPpwwWIDTc
lItPpIx+KZB+nHsEUwLTu69z/rLXitL7NzWblLatjCFIfSQUVigORiF/w9U2fmLCN3MlZpsf29a+
v0p3l0hWP9jGEZndo8EO3Twksw9v2MZHzoCwWWIXB2hFhcNKBR57VpXUWD9DhwG8RQBv+FFVMoyd
FQ5Qhhdm9Plzr/ucN6lwiXWp5sqekxFhMnM3RMOX/uuGWz7cXa6wVzadc/XMhuabk6sxvGCpmDgK
pax8Utmtsg/3C7xTcsXb7/m1utBAfy8L+iQkS6p+vK6h0Zo7Jr3VuM8hPBc/Z/25cpAxgXlAllEU
JA/WqKh3kxMWF9D7kP5wqdyB3OrEoGlVpCzenoUkSthtVAqq82EToMNm/58P1t3TlfYaq322svXH
CJAr7mV2oa6nBAA9dgJiEgPjgo21SprRVZXmdSpggXgOrqbiTe7jPTEajrAszhKTA35y6raLGRw2
z3ig/9efw6+GMh9AnWiXyMWcLfb2ipGsgi+6Rdgk8T9GI2Xb6PDqGEdnClcu5Aq1SqOeYhbjrY2E
NsNdYsV+GjPYzarmOYfNTNhULOjMD/9U2aXso9u34I1O2qnicSLPJclw9xDw+hbBWTtndxu2SLLs
P0KZPAUsfAVwSXXHnJKaW6XP7zA5e4kXWTGBv6OUR7rOgCyfqYvIIZal+DkjCXQHiE7e9u8Vuck3
mNYhANZvFARxziPdR7AoNQHXe6bMDaGG1tEYyGXk5APLKXp98zTSLcuIN4Rxyfi7Zh4Q78slXDs6
2dKuDBch1NaFHduSvylyXJeRFonVhg40umH6YWjsSTtJC/zERy+PRrZLU/Gp0UF7LUqUfrcwcmvq
Brtl0TB/75RYK23CExm8Ffs46YmouZ/enAVPzdMWgkBmUqu90xBDlaleDSaj4o9qQESS0MOOXtBJ
eUU4ikBtkMl8kdfKzCd13iLRPFznFPHprp6UPm4bfhWV1XR9IEuzftGGO9H8qULBEF7PTUrbO5Yc
YTfY9mATTkBH5Gv7tBY0VeNme4gF/CE0Uggf63aoEgA+LVUzRcsqvPfZ6CdxfbyuKqUJJ2PuA7XO
GMPU0HhBpNsZoAc/rObBzPFClaX0MeHTSC9YO2bX/2suUZCTl66hLpS7dPUaI8RNO5sq6jYQRDqL
Vf/ahYxMkOkpuzhmoMqJV6GcmAIsmG68HDYApbTcf3Nym9k8YUpgdd4cwJo8gN2XZ/qp21/2/rZ4
pIl7n1LC37MlQvmJqdZyA1Sjuogsgk8EDpURe9PdWrZnJypbsTeMNm0qZ4N3u41EHQQfGU21hcIe
MvjBMCCzVHrZ3bltru6uqcCTgkDjYcg4B8NfhWkdKh5ywoZQCsg4EsPFTPvtMfSvC1NoOYaZVufQ
QW2S6I/A27XMR6OA9dnLBibgG4q94FdRRwBWq4g45IEQfCtnW4WZ+cfWbpLzbBkyghsvWGSJjm1Y
A56uawiuhTJALjMxOULVjDg22E5Y62ZH8Kt2aE0erAW6just1o9F5nKJUps6LxzXEcH6splSDN5o
N2ix81ajU4SeIB+j2tkSHXhK8wv118XrsYc7xsQYstAlrVXNvXpr7lgoZ8vg5E0hlShhx1ZXz9Ed
q+RFfykcGzh5Wf3FvTLLRgmYYfGfEZLJf5Q0e7bmZJ1evz6LbpSzfeGvreVipkV7TIkfMd0U68H6
IcgjY3ZkT5VRFqDIusfD8dTEbjcFZOK+sD+u0KsfsncEFAj4orx1BHnjs3w+txy62mRjY/JZRzbN
fxMPEeZQeaZCmwwvPgVawFh/+2rIw8HBKQpdIA8pj618gyKAj2a7IRJixuVqtrKZ2GxTaVXkyhTC
KG9Xtk+4XxbopH7AAHb4JNxxgEguDsX6FbQM1wfHiQe/JV290Y72RrFbkS2qLzZd6zsnRAXoOTKr
5vRSiPMBVCiR+na/y0I123j7Lozyn47kwufMKM0lThc06btfWJ7P8Qiabb5In8IoLRbsinGNr1aK
4rICVpXkKeO4zxRT9sRaVD7Pk20eFUkCLo0NJfGbTMA7fy6WXmq4CLlvHHkQw/JEHAdK01W6x9vb
uXOQGLoYtnOCN3kzZgrDDFF0b9CDtXfj9kVjfrhh+kT2PaAdoeD0Tu8MmeXFWbN98/R/8FCs9vT2
Mxq+iQDthN5E+gxryveIZR9K9s29XEQMMuyO/gnveaf9ZiaZ463Nuetq5yMCy84U8gNyxEykdGGQ
dECXOuS1f/5Kew+nlCX3TchU1l7DJp5PnW0/F7glKAcv0EYuESfVG+e+NUO3g774ABzBpv/SBqAD
KSpi1L6Q9LvDX4O2wF+a18y2XaGhHx5OkNbRLJB9GpI85lfr8TKXx+MvWhNeuv+NxI/bDy9WDf4r
hn9xPOBdJa5gq0yDdhyvkU8ex3TmbOyDBFZ2rI0ixrg0w1G1ajdJHfBv6IQwUzkSWu4+3ROBTlxU
9yizZWIY8yk3ELv8x6tqEJAhtADo+kqcwNcJX4p+hiY607XU5fTBO7dP9GqTlM3cmp3ZpcBXSG4i
/mDZhd/xjN20trp7OtUXLCSJSL0+a8Zlcbfv081Qet5BOnQ01X1wcNPqDt9n80kBq7t3jfJxzoT/
ORC2+e44V8JEMI1uLtcyB8eiPKUislgp31mb9S8vaFpTM64602Mh4R1r8qZPkU019DRZ/bHEf/gx
7bHmQrfAS4e62peQW9PPsLO/FARECjNvxEcrbGGo6ut7KgmH2MS3AAwHOTBtyDNxyrZmJoAscNkp
kiaxFRjfPBRPtuqUEvdvEVnkq/IVgtox5EdFXu9zRJN9vsDEOz0M5wOcN10ko+KaOu1vAMVJoe6f
PuVlzEz0QhaFVvSWiyhYFeqRc6b9AblokdQiPtRi9Y3gH5j47cLa8+d15qjdJqW2YK4PVDYYqJQW
tOfzY3wU5bSm8qxh8i7zI25Hm+nhGpMApDP8G00wfZjYYaAJFnyOnJpJdI293nvuk4y+LRAgnky8
rDLonjgdridLJkAi/Vd5IgcI+a2GtxzVjhF6oI8sGNFAvTAC4HZThWZMc83PyWcEUtolc21/bJNW
gW4E+g/BkfAo5t1sPv63RvD4SFIGrn+IcM1BIfhSDAWTGtclAxV13sdiv1qQqltSIA1LoVWvLXM2
UuH7fWb4uAF7UAZ10nTPdeCmzdYgiZouRRpnlV5T8Y4pNxo4Z4KOefevjSUYzD4LotmUEAi34mFc
xTOQ+BpQxZprrp6tBIa8AzTYhQLYBQVeb1GYjvehD/ZmXLOfK55EefbiTj7GRCtkAPRI07VJcUYD
dmpIsahlKKA4vcL2ZX0s+FWQv3TxWX3U5KxI2JmBe3qDqoz94rSkyL8q6owUv95FwwJA7QbaqUtn
P/7rjMoOsBY4Q2vyK2AxNlk3JEgbWzZFBE03rIScLN+ChfN53j9Y+srZhP7o55GkmGJbZUAc1jFm
bgCRpBh8CQKjcZZpNLCIudGEDICMzs/1fnOGPm+hGK10DyeQ7Vc/UbR29lBfs0rfYdJYophAkCnd
k6qGmTzUVumuPkyun9iU6xVrOGasX/53lCNX1BG1QDQCaWi7+xki1x7HuokALYB39Aeqj41VJqBg
wy44FZP+lcY0fZNZvQ9X6uPrQDGBgHoHX+fec5PnILTVFHpIFgngVLCPWtoAcR+tNP3mO37wbhkD
0wgaL4L52i21JS+IMj5cnKwAxiNUez1QzqmA3Kw8BoT19Kilnp39TaJBxr5bFTW5nUuHM8w82542
VZZnkJA4WZTVCdR/ExlcrEqLarZ0N5d4JU80X1Ok0cBpanH17uZZssbJCHRE94fn8xhrkFHwMvzR
EWiksjApKjrb6dQcs13PLQ7WgcscVyvQQXNjHzsHiEy6NxWPt58BMx2i32u8vfvdUHU/KRoz168u
Y/DkmPUZuYCiwabxZT5yHvegahPmin8y0iR93myLuCAx0je8fqNP7l1hm71umzJ4UpTyASJyb/f2
DTXcIRwa+UyB0PPlHDdriR2Rsb1H5oJwbGc4gomqLQb6PLTPiSwQWKeB3tW+lq4ig+aKdREjfpww
PW4no8PBDlrZ+7rbI33ERIQbKdAoQI4AA52avASMCUZ7Gtp5URJU4YEyAWfmPFqeID4x0dWDzljZ
/LymAb+bJnk2pJdaBkDEsigThsYus+RQRnpyw1xw/eJNy1mQQF0WkCzO5dCyZ+reQ1PcNkq8Bpx8
smILGZWkPS0p9dRWkt3rviXvj5cpswa1vqsY8DED8dQWfwqiRrUhE7qAMdPoR8OWViFVvP9hz0Wh
la890iMV2r/YvHfymbfzvVV3GG2+lrinyQGeSftQBiJn/Pjx8ur2r18bshRsRJy/k9p5t8oJPfok
dBa3BcnjnzXlZg4hIb+O1Utz9kH3u5fiupedpFHLwL110EwuAi+Wb06Xv9qarZzvR82MJ7NdsZOm
cVgoxeONLENmSLlf+BRnQvWd96NKbpGs5rQfh2XpIb3wIIzEfPGs3/ePb44GbJQBoq8BxQzeIboD
rPJILyI3IARoNrsq9w2dJunAGhDV6tTQ180Ct55jbspq5w1TzOq7uwucsRVM8DBmV/2SZ4zDU5xd
8OD9k5a6EBXBLAz3L/jqLcU7xUCiwRtnB6qp9slNbMagTz/1GFr4FmTlYJlnlyUIfnkh/ajihnni
YeWE8TiGY/rBQGg5r3DKQhvKSbvybWcQivTQidJwdgth4qYWXK7MKuDgqkPpqoWVODBo3na05C3k
PIrVJyssvAZ/6QNW5jx/04Qv9gWQ426RmD+52WU6icXc3m8o+cxCMEi9mw/HEndLAZsDopwaL0Sz
2mdyRzqaHd7Re7Z1CInzP3lKHoZ28WU5VYs5iThWm5tP6UxHqNSXqaBhXmvFuDjLVzlbXwm+d7Nz
SQ/FgMDbAezEa8yfbHok5EJJue/c+HmyBxCGllswUUyw3b7dJqy+AT5EGAhvuT6VrS0h14jMnul+
h8bxecMkuv1u8VYcroBVfpAO8e630g8QU2v9Tw+qDcWvigh1LqwhmgjN9o4hSORZZ9seJTP0Y+kW
7CEI0Up76dzHLdbdsbEeA7nkHSaf6uFVLGdQpGtoazNvpFE/TMhqyzlpqnLWwbvBt1ewyAxzTXMW
OqTIINafL7ljN/LAPdgGSfcnUxhvU08ErC1lr1yGrK0aVfeWznJUTnEE/zT4SSRyJdFRpIRyoN99
Mi0A7Be2PZiV6ukgCxq+F9wsjLVS5Yz3XykO01Fsn6Ng/DU0J8EE3Xc103HG3fVzKqZMC0KyZqGf
G0sxSdeYl0pQGfUw2XAfOFHnybwkB99WqodCTrWo5gMneKdLj9u/k79rg4v5Ge0NY1CC3uuN6psX
AEj5Qbl3BEp1jFbJnG+YmB/QLtuVGndcFW4pgHGLBXHvTGRkpP5sAW/hJVgTV1Ixa3QAXcTkdbIw
PxnaasAxd2M/koynVkArQjF3QwFK/k7rqeWrFCwL2P1oQeDdJVLZYw5f6rUF2+7y0zsZEnrVVfvo
U9G3WPk/JzVu0msYdPw7a24DqqkhKIAPjNQlXdTIdP3+6lU3iyiDdMlvXEl/u/NF3EwY/nZupSoD
VzRnzTP6HpKU0/KoSbH6EK8M4Ub5F5QMFsoXMKD8X9oVm6Nxoxz6RHJw1364DR1wyNLzZYvXB+HZ
tC/ADCjhkhUlwO6LgN2cRNSj4xVqcVhCLWUPBMZR3CFBMBZc0Tc/umD1dEPHxt/a85+SEg1+nwXE
ey/MT+SuDwGc7WVVrjI94RopNDFbOpSEtj42V/Qd3j+8/mCB9BveoAlIXsBtN2qKltQmZ+3CGZog
XOiqmvrLwomDei/hfh3+EsQHW1obS3fapiVL4ZXvNMVNyXH7aFk/z+hqgh7BJK270xfdrwcl5izn
DtCMDf0XnlDwHOGao24BAF66usaG5EqlXgRm8lbwxtMbIwBK42Dne1yGVfeDVYqyfr2ORdRmScKV
OcX6b5pI0Zmm3cVdglxMuz9SYe9+SOxDs7JN6bP8y5wv4wA3o9ZHAROD+LOIDtYOkV5pJf64mQ4W
BaRq1aeYxTa067Hr2ZkDFZ8UFNg8e7zeQUl3LqSTOtvcw97i7nLI2gy7AeY+rdU5mCdOLCxGpxPQ
2OI53crE/aiMVzRit53nfXpYid4a8H8Dzy2o2bb8BOvIt1B4G4z6aOiPAsWdKLhQxoQ9TukWGvTQ
XHqMibr7GDDdWvhL7BvClD9SfY936L00EUOuXOmFfElvsOI2vlhJBQkAboacrt1WWms6TU9WQWYY
sUB1qTPz+bTMCBhj44TfYHPgz8KWGj+PD1ykb88tmcnU0UGf92Cwo8MkB+I0SAljXHKdALu9sYvt
RcU/9XZYrm6Ib2IN2teW2Vddm3LhMJHID0kmO1uus40Sq4pkOjAmvzSlWm3hYnwOJcLPw0YRQoxo
hQAGHmHGsRcthpWcqj30GLu6H4EFYzoxZzf+ILDr+IToiVLN3YGlG0V4aBsCgmS32qnRG+Y/+XzW
yBgQVtu9HXUfetblLnNxNHyqA3NSwc0NHcliE0NbRz6hIgnquGiApNi1l4iPPobvpu+VxQ4Vz23b
+4clpULuHSH3rBt+RN/MiwlEHbLwsd0XFW2uWzJekZzlV1oLOP/7/E8cw4ZUUX+sSo6QOf1NH/td
RpPEL7xaD+XNv1UrILwLP7505TfXDZIF/SlvKxfMtpKTyGYhD1HXbd06JqoWoe83FnYqaqD68sKw
T90iqMuEcO59lEFQiNeqxp6UYhO23Q/3Ve8/Kam/oT1bg6GPeGd2hTYmTJO/M93lYzznVMKVuZhQ
L3qOiG7CjV38qeV3lJOKzG5Qpk5je7on1GRUSUlUcdOqvsTRMB3Y63foCtgwPawswAHnK2kX3Tci
JHB5tAo3sCyylMqGHWStxYlaVz65VPsLosXqWejuKPOu6T1ZTaRa6vnG24HQO+NJ40c7ewBQEn4B
7yIWf0YIYpHb+/6Ea2eAuAP9LPX8S3mkHfPd26/nqpi6Nzcuk48rtsVjYPdlf7zZkuRxlkbNZDRC
4yhU3lH1VJBs0fR+93FCqEakEFmaYlv4D0sKXMhgq7USFEuuZBp6NdY42UDw6Kh5f7CWYpl90WZE
Ifx/z95tRWmRLie5risNs1ExcAJNnB8rx/EcB2SyivILO0LsWNDY1DIh9kfflZ4BW7ngW5PtmzzI
BWMEf7d6JA0287LcjZaanCJ2swucCl7SyEOPtSVET+Xfe9nVJZu1l0aoKb5gfg7oqbf8m9lPtAjS
nB3bPwkjoNvxgQkNvCtzOTQoi8oszpZimRCvLbDepYQH6FV/SCYCscBq1D4KUzVDbWJH0enxYsJe
Qwi8J3diAW/HhrS3AtXZtxYRS+BBIO+CgDowwFXNw65YPfdYM8ph8BoLsUKac0g1XQ9dDJxor0XD
XJKAuzTbgYa6Qdk+XeHksCXLlG5glT91UmnF/PoZpqTkkV/ZeCcDKLgMa6YRn/Mn0ks+gp6AaLlv
ANHrRvxSILoVcZ41t99U4yEMNikUHuWLZklG2GjpYTgII2q5uhwFeF6NQstlF28yX0WxGuWosGxB
4j8fJrsFdROO7oHgk1ZsuJUOLfAdZe+sHwpCDn6uEUgT9xSh9QXeVVUPjqb225fnreHDyaDoxTnA
1MjmYA5wk5Y9aLSS+e/HqaJdtf1Z1SCz6ZoeC6nHrcsN0mZmhPPkxoAOO8H2amcRIZI26wiRorFp
S8VLiBknkpySnX7v/M8KQ2Ju8ycEv0lAKSAoyZLnzeu6nElWg74BKLbgOvhcdynBaex1vdOl5Hs2
IeRi8IRUc7MslsyFk2QHJUjKh8M577/biyjyGlYMRKEEy0+BlYnLzqSNo/LEAauEC6lbeMRZJ/pS
o0rsYVMLgGKGEW5QZOFbW3C4M3IdbUScH5LdEZJU7sm718qrvLK+o7lb/NubmBDjeL6kKADY/mm4
9fU/CopBTswmacIHhPKF/QwKyx9h23j9RG40hXHmZMXssSCUOO1Fh+xjvV8fmMlJ8uVQQvhFbrk/
sBxPJzyjF8PNjr6PN1S7xu4yxuQ0oK6Ky0G2I8U6pSZk8q95stzft+aAfL3EY0ih8v+Ijc0MDKlB
QuM2/yx5XloPKZvO8yDiHnbcTY3TbD36qiTyA8w+8/9MZzYov3egwHakKCEfzm8k138AMLTy0ChZ
+MjJXI43Ex3LA963vMtoRTpNHejQBw9jwuu4DpCjwYtg10Mb1DwYMDHhIVtlzB87sqFVpxguEAa3
hHErs06R7YYX1temtwjKySWDpWx0AUIuOEfFE3jZeHYFUCippojcelzf0Ic/0jNQVd08LDopXZ6D
HzwOIXgggXjqmjn6n+C0HrsjDlfYWNWLDuMshmyKtbhzA/pW1sw+v/35hzXBNOUulIysFzXYACYO
nRJdCcL+gyNKKVhfqyGZ24uo5ePzoXqhqW4u5Wx0dGUSKC+Pn2DXSl3LD0AXlSC10DW6vak7VGe3
aZLj4l7X+ml/ixgGQow2JgNNC05OZiYvT51nYLJQWLLH5L/uHfE7EYsxQ/TemIzKm8olSO/ScVY7
WsWgmnryRUDgpoKCKyiAYpfq4XRkzK/CP6jU5GsfPRs3SWnHay8NEvo24p2cgoOyh/hBkqege2DA
Kd9jWhoaUHJjBl0mJ5TneMYRxpeQjrjG4+1xQrQyjLrN43Tec+xzkjYnU41XhzU1BZCxQ1Ziiazw
Bt6EVM8276Z2LLGDqo6u4ZHCWef22V5Qqfm1li+rYBSbvKbXUE7DSk8nbwovWjH3jatShwodqcjO
Jz/Cud2bwxuKdmPNuYVcZwG/0idmGkQ2Uj8IwJ5y0LU11wthpSsMA2zrxiXQB4MrCWVU0wvCN8Bf
quNY0oHgNCB8bZbxshv4Of7HS7zAKFK0KoYfLSvrwv0728XuvjfaZB9BKNJRLMYzYmJMppopW2Vi
MdmMLRcRWkmGpQpL2FjYywGu/5BXuzEei5muA1ULG2K9XkmALiKHXX1xusSGTQUZX0FlOq5mwIPL
VA2OqfIapPnh4r6cPM6nbJW20GftW8xkDHxaYFty5LuA2EbWV08gpla9zAw6+ZFIJuI2XCtMYufn
Nm1LlA50xYvJ2Pp/uxXJFa3X+uaUmgpLU3mvD4BkVoocStpV3gCLF5PvvVCE21/iEMnrXPKOU02b
32oH0qO0lqc1gND/Cjbj/JEAzFAJCmjkrN5pjRxNt0z6SXjdEG1iy1B3FOYl4SJZMsC67fxUEmgE
fq/wO5n3N94dsSJKUUXak1G83djZPGy6amfFywf4/VD9uEi7q7RdqeZp9VuEp9xtF5APIXXgp2DL
ZcMyFykElDsefXgosO4E2nE1xqn25aE9kilaV1p6S8tcmOTXbeZ328RqZrohlMV1/4Qz2gryjHRf
QAmBiA6N0LVwxyuu2JYwnY0HOcu8zsGPEer07pHvNHtsG8vfL5++AkFpsSrrjFnBnYgr7y01yf6E
bNNOvO8E7GZban+Xw3ACSH7HV7qSQvxRAX8PzxuGim/8SSI2ljzmlv0rhQHOdT5vsZdAFIwXZArd
IAhwMFswWJrDjuINzUsQexPBWFMAyMs8rTTuaKOiBr30dHYZgeKYOE3MUsMmql7KeOM1YgqUVdf3
yk3lqikWJQTJhs+/SLF+L+jbwaeOnYic6vVfzl4z8n181U5IFNHA54ug+OzqT3Btdv1vNb5z9FzN
i/04A2SbHIDolM+6KpuYTtBXpQ0wRlMrwCwCfR3JSJPJUSs/wK242QrnTKDgaFl/duCHd8+f+fxI
JwhpvxKq02JCErxfBVaio77QjdOr7EIUDl/2IzkC5XkvQK7wL7DN2hMwpKg3ukVlx2G5FW8cleMG
FBCh69XMJyBRfs1owptcBuNt0dpWTesaew28eAUh5Se6nVZRfSyNOCbUnOQZEQkDNQiZk8rwEaU1
G5HyqPvagdWSCtWotc8jtPgn/gymgMaA9gA0Q1RbakR8ZszxucvsVs+3+XMKs0IspxHjrWt80jei
s4etmK73YPnrROQNJzewvmpdlN/A3Y9WdyD6Kzd6sRI7e0qq63Na4yHGQh4RK/XdBqPgWSUcg5jX
9DcEjsbCN4UBPXMkwAqPXU7/IMy7Hn+ILTBYZgyKZRtaWCbb1cQoocMwLIqrgWkcXNbZmK1oAZrK
YrFVj0Cc90/72fiVUuAVqTc3YzkmTNL2bI3VeGaF3jbFvu2uEUsgNEtWrguymjPYIStaEg3osLP6
qa0ZAQvcyayqM01JdTxbDCLqO/GE7uCGabUO52A/lZmmJGe9yDXB6WB5ImAh43FO5KyGjZBZlsjK
L8/7NAuyB1QI8TAvsnsTXkr4yYoSC4Z/I48pgi8DurWvEHyU3hMsaJ40RLym6WHJOusyFCejOJxv
KOHBZRjI97oOaQPkRJsHfA2J9nuj0r2SqIUd3lnTZMeeu585yl1JO4rU990UaYis34T3wccHCVDZ
YE3HRapu7eS4aatbwERn6NCekXBN//FJyXRQ+7jMRX7s4kinIUD3/3bBhWzdNk4XpoS4zKQJccup
7YnlD2fTbedEsZDWESL7T5nzwfp4JmENasMVTsM+OIg3v4LxC/gUbb4SKFz/Zft40lTTwhPStN/b
oy7T2iEhOF4LDfi7unEXz3gEpOm96uX+suR/bsLGxgAtb3WR4Y+3pNatR81cfubqudumEk3JD873
FwdjE4C/pwNxpy2DJ0hwqPVZL00tY+JzZtvp884+B5tfmF8J8x1vuqLAQTz/CHEXHaTqI+v6piMn
aevGY4GwzPbubOsG4NxjqV1lCplgxjsHpbVXjWAV7Y4ezq2qKchfBK4BfG+8xJPAUGOTLyGnZStl
FSldJV3AbJER/bgK0xWCMl5kVrLgsf9UOZJdjeFHxILNXY+tIkyVwCIre58eIV2h3hpPoakNdTyR
17MqyLVoEJ3FFdWCemZ0TMF93iDOamxf8Hvj+ZEveaNZAiymYrVKtsgDKmTDdHNyWbE+Tupb0Tkk
VPongvvbd9gXmO99c6gER+3mGfFNNODZZX54rrVL+FCWo0A1B/0KIxFd9eiJNmc61FjjREtm+cWD
lUCoxJt/w6iyOalhGQ/qTBwsorHP2yUhrzQ3Re+XdHM5sBPLQOQCZT2llp/RkXrd7zIVgz/qikMZ
Fs7ABBxKsMqZD8FRO4kVPBXuWrf4h630tUMuH7LhZEMHn00+7O04BpSp5Zc/Gn8ri6rwbmEMfKVx
Eg09zbH4I6tGKced9dR8JZmII/xXi4ytnrdW58EKC5R0fn5cvsyf4SXlBCRKdAtbAc1TkC4Ey4nU
7+ohziNtsguBV+r0h11HjQn7qOh2U/wNgJxwBzNH4dCHTC/rDDV3t/s31oWTHti10nqVtsbmGkzT
wa20lLXpeA5XncEAqSEV4+GpLw7SyqeyN4yav0AzCwWszvt56sd2pqjRvu8mecXT3d2vm4ceDUWK
Qi3BUkrQWIaS8toIkbuFMqpFjiR2tbEkKYSqc7hmOWN5jvnVMJTUJZ95A19ZPpf6wZckNFOtvayh
dYGqxIYaB7ktOSrum/uuUVY33SkWDSWjDgpEXYxE4NBvsKbKJxvY1tpAzOgfe9cB3AIiyPA309HE
HGWXCSPCmf/tOFFT+aigkk1JPZ1e9vBocTwP6LC8Aq3QlFrnAoblygvXu4ub5RSNp/SiAC8HMcve
/8j5GzabpAaEXMqXzL2RKTzsIQ6sc3Ub7xYruC+TzMAlqN3z3CYr+ErrWohblo/MNZOWJ7HERm60
t0trYrBehP+xgS6rty7Ve0v5boOu/YXJ314U5o7UUlcbs+Zpx6ihmbdtfeuO/6CBQ3FHCDIwM3zY
KS9tGk1sgtgCrvohjasEpcZooN4BRvhlmfbozuHer7x45AfLL2BWfzIJ8JriZthO1e2q1p2brR27
0et2kP45afQKk32ZTfv4gxPUwR4Ta3FCtZmySybbHRtXxbnxvnVpgwApv0cFcJAoZk+Tco4/yy8a
sAFOWJMTu0zCnz4UixtAzto1QDzxaoezQP3Fp5Wnlo7rALqBwTxl0zmmzvruNjlhDFHPPwTWkItM
8b3Lodi+iRhujtdk3eNgJDA1dQwYwd6PT3VX+LkXoW+gOGetHETGEzQ0O2Sa8+cwmde7htAcRkjb
coEkIcMVW0RxL0PAUiYwayJpRE7yzveJ/GDEUyPlI9oxI/e5DXeq0SrPL/eAToMp6mfEujKSht8r
fdu/pYsqpay/0vkBkX0WEjjQ0bZY805u/mlOQbQcOvUy6C1AScA56D8yQzNb2yUCodBt8bIOWTIQ
dlyr3SdICzZ88FBynfjieSTdpGl76S8+hxtsl3PnbX+moQgtIMCv83WODjib30lOruDyl83ZbYEz
+lEloKrQ8sh9SFD+weuOB8cd8hLhlAItepl+x8th1DkyU+I1jZMHACKFEwAN9+jXKFg+A6O99rSp
AWsUxvEtcwp+oG8VL3ojX665wZ/AAllt87zZRhcXqlpXkcy0qZTm1FdQMRUWH43cdnE1hViaR6A1
iNW5JbEe51WrwuCTiQ5fn4FaNm7xIuOzVD+c9yYN/228Xbapvi0VU/brc6y2ZILge8pJX7tj7Ip5
801V8pLkRh08tIkln5FJadI9cPycfXEPdONgQFQJrQmOJj7yCpxFJ1EC2NIlVMMLbN0Hv9wqteI9
lpzlHUcYmJ9G3On9RKmJIkwggg7j/mW1/3y8EYrpL2m0lEQ5vZDTm83bvQOwLOKBZvvRRRGvdP4k
IyqwokKMpoHD48IfOaBpFqijV/04K+bT5hJ7OoyNbER9D7HmMoKzCpoafuTc/bg7QiZueRQmwZIW
J+mng35Ht1re1tS4s+NpgOccmNiB+2Q+iPg7MPOf4bVtCcNrMpjugp+98s0WBjl5joKK8zyS2o3W
Br26zkrzy0zJa9KvJPGrFel1eqs2XP1n2bTnas/pKwNL+v7OcfRSN0bKuOmaDDO5gA7cNl2F/pim
mnolk4LZUZn1w/Fo/YRASOU74pO6HVAO4Eq3u+RmqNqFKUtbosEmRyMR1hbTfRLmslC6RaT4N+J4
pmFVW8xs82Ls8Wflf+fxfu6rIZKP8Q+H3u0e0qEUE2gIV8Eu3ZxFVw6ozvQrU6N+Uc9A8Sf//cw7
2qtbz7ilU4Yv4vbhhF/gXgCFI3wtIe3243j4TojVepaMgWXMKE3Uovi0rVPgL1jDFvQbi7yFUHfm
yMe5aj5C5SOrYUv+b3TlXOKzIKOXF/L+uulMTu7/F6WzchBiI+4O5plYEu9NEhIrV/uo5zNfMl0d
0l30PTfp7TOPz5iTR80pGK3fe85aqYObzpOn/m9tCeq3f1moU8EJN4dWKtc58qxs1ST86rBGk75l
P/a2TJjY+1g4pBQw2jRnuzY2+5+yXQe03/iqA/U6uKa9Zb4o8qb4GKNEjnPrZ8n3RsSzB8J93Civ
xWN4zU5CLe37RPegio7FZOY9MV0oO+MCCHW/6fPJsWQkpFt6o+RfmjWvPLJGssdGqtJwcE0U9Vii
Aq7murdvZ6p46I0h7jPgyCc9faMW4oXifIXz7zqkdBH8Da+ntsiUXZbN+TZ8AL4O8R7EvgMos7VO
GdQv2VHTv1+/Qt/LtJY/Rnqgb7PvWkTYevvVuObEtdLGt6DZQJmcY1AWcqTGjzmtTjzrDz0aKpCA
r3sGmnvZvWubMzWGLX5RwgMUse3AtojY/qjvKglI2+IzcNOmJBVjoIx0sQmNeIKDntkXbCv/XUF7
U0QL5CANUaGZvgQrKaOrNiCVitp4pwKG9Ot1jpeLFZs1ivfB3+XxEN/a5c0aqpSf1fzX1Fd8ktEB
xfOy3ir+merElt7ZYK3TqXwSEq7kEaj9g9t2KP8WsuemO24LxIY3+nVvFro5DGIMk9K7phiWKnZ3
jl2vhKRRMck77wIfKVmUUsFEt6GZeLOpOtBccFfO2wgawH59dqR3j7K3VerJGNm36Y0DeaEu8vYg
0LtTfw9U8SnJ1QWuIg4Pc4P3gHSz4eqgtqSUAjk/5VuRTPlvb3fK7LMnwAdRkO8hrcyCXCPvFhjv
e5iXX8v2PU7gpvTEja3dByhLKCMfdx07en9MbL2tp/P+zZ1I0QkVCgQEEx6li8fL7h8LP5fX+1rE
0WjFUpZEfb3C317hflnVmcC0pMvIyt32N4zjDkbqte1oJbQ2flzM9pzASJU0g66Mj7yV9joN/Vp6
eVEMpKXPzxQF020i41ALC/QOBuGwpeIIYKfYI2Mjpbqmu1pfK2HG4KNvnSIMIdIZ7FK6TncpqRIT
j8bz73KvkyMWC3XcgDEttmE9WN+eA9hpLe6zCAmMcKSP3F0q1sJEv/JGBfd971eeauGsD/cNrfE2
2NOpB+E/74TEDQ62UpKKTnjdwC8MQaAQD0Zj0PFJpnyTlrojxRwiVi8QsQqOVJ2Qthdy5hTfNJdp
pE4vfA2R/rjRC/4yuCV+IrPIWknL4yY/QnqvZUndhj+xJcpp2rCAX71q9fstW5XCNOnOHqxLzUvF
XfpBbgHohzvaEsBJUzqUfcxJU1cmvoMRgY+ZwONPNsfVWo5dkq0CaNGJ607wEK0wZrNHEOiu0nPs
MJN8gJPnQDQRM+Z2Lght3tk384uhm5w9Yu2IJVJPwojm8bQVnMGA3SyoKlyMeN+HqO9aUhYxZGdH
qqqMDSzI5rHW2YUdKJCLroKQut4tE1P1wSs45Iziypxt294F87y2x+giovjDuDjp0m41GinwAm1w
Poke8cTCLjk94nas13j2rtGVMo7SdFAz9NC2mmtX/vzukpviG3jgSGSJZiNJdMNDLcuUYugQHX/T
ji+JCRqtQnLQaA72H0mHyiiCxGLKK/3748zae743TlNJSux000ABtkQdlrH4HbfwJUVACoFkA2mA
VW6NKf5SauEq1k7yk5nB0QEToTbD5UagMphKLLtrzDY1Jf5tZQZFspFG1DOJNk2j9fZZ3GRUvqBg
gyl/WfDlvsSfJ46KbP3fESjDYVFWIe6y4j5LCfi9QfG1WBRXR/cCUUiJ2YM0QhUc65s/SOVF2fPn
NlauX1exFTOky0B/hsPca7DrLWPCifHgco9yIeIKM4kLAm7102FpttYP6IIZZhX0JP95FkMgxk9V
GHPKRFD2QulmvsfdcsvoiML1npUSCUA+pNe0VOv+TV8RAcXk/V71lPcsQqYANTsIujmEI/CAbm1P
5cz1tlhjE4RosHj8InCKu1gF41xi7xeF7S3VhCF91bfF4FUMeOIsoCvQZn9nd6fRZQ27vZdllhDK
ZQfyG4URypUXW5h6rVdahiZpi3UrhfW2LBNw0l8q8eCINPAg7gEQ6eBnp+vCjP6USB3MW94ltDPK
DdHaMHg749igy9Pr4MxMfIrej3nZ3l8F3gs9JL1YLDeqXJUt+7dxkKcx3+QKDbvX4aF35mtzFFP4
ovRDoaUGYoSY8l1JGWhi0zQB5D+yNqsWArM6OoiCM8Mb7ll7cBVYtjhvzmQr2iVAL/5nKlU0/kkT
JlTGflelEEYt28yFsy7IgVHt+OCUUelNfqo3hldKyrXo3TTC+uVBPB1qprCMeMMKehRlsmaoHnj6
1g+XTuIzDRqQaC3AT/AB+Xs4tk+JGIrRIvbiY7RVmtSxbkIOzU6x0mSRBtEylTXn62mFRarLj13l
MTYMSRq0lp9RmyqYeVIKAb5uOvDkVL/q4xGK/6CVTdMPoAPifeVeESUNkw3Mff5/cy33/kZGAM/d
zWjLAbivJ1+ZwxMdcvRUt1zZlSiatVUx9qewpRenyaFkrli355OapITAqIiK0QDkUxFRQe9jX7Ig
EtYViyuSHiqmYzTpjDbQcNJ4UdgW7naZ9GFAPlIhixZE9DDC/MYHYI5XAlokYQUddN5JIjD7txvC
LMTYjI5r9sI33PC4LNcjYZNgRVaUbNPnbX07H+mNFQXgPn7PYd+eTeMRoZgjBd5RodqbM0fNiLTS
AwOf13uxQ2nrVZPdo5xb+tpvkcvyY/m6x+CDBWKFNVCEd9ns96WbuTb0/ZWEQkucdd7axb2yMpLo
868aIMOR+9+0xUryd1QO/ndyFtUj6L+EItahGDQVHaeLOz0794jo5sYCwKCJO9gDwJsmJqKjzsmU
2vZ46OilPBmFflFGihAZhSjx8CX7wP3JSWCHmvqr6JFCR18BX0RJGMXqEfJfBJ6ngP2D+tl2eqBk
bBbqB7hEwtqjROAMBUmMdpTdCoj6vbyebmssSB64NO1RBbiuEhc5PZy2/iMSeRT1yM8uJGF5W8t8
sveYErl6+WiLVS8QyWzXrzASq+AU+PN4nak+fjIhDvbV4cH8/nGRsT+V9Osvw9Boht77JVsE8RnO
WwkPS68uVG1tEExX6akqhL3NiFn+oMS0LAKobS7TDpQIAWpMXscRNrDx+9E8KVny5AX3RZYN4dKE
xQZADmJWu1jzDSsl+a9ZVM87hGXWa6dlDRrLtTATLWtKaKppPSC6TqxlmdTVH5OmhUYZJjm9Q4nq
FLfECJ0atQmWGUeYoJL1pkh4SrqcXmVnD+MnXK3F5Ot8tFI1Q3Y4NXSsEfYvIIuzbUQ+xHSjptom
+Fz0MiEjwoO4P08Mlk/r5xEsmiX22nglI/OA6xbqR5fuBvz+GtqDQt4nyyD4pHBSNrerQjlflz+U
EK6+sdXGK2qSdHWfrH8gHxl4EK00dronZBICA5krb4f3IRY5Fp3yZC0nx3YJk2lxb9g6VInTmJ9f
zJ7xiScdg7W6If4h4+UWIZ/EVDdKtJKKHWaGTc/LC0KtAKZCqxg7y88IdV6BI5PwrXF5SOwzefPn
2QC+Psp3xsvGoQDuaO8qkyfWUsy5kQaI7x/uZg3BVMsTgrwPJ9ApL8u+1mMS7aAKiur3v7JPD1yx
EXq/n/D7Xx2H2tI6v1K6ZisXrbFiOQvFGQOV0yayxT4d8nR+Bzk3rlTsc4n7ZxFfqLt4QR94/SIf
Po6ML5rczIkjpAwW51nqmElROhblpmfC9F9730FQmsd43AC9LaNEa8Ez6BrFrkyN6WkfKMQSE94b
IzReAI+zox4xGONs3aRRWhsQPRrHFA7MtZxnMSLHpgNcovFX1hEPQNhGHqoq0H/+OKekfK83km+k
FqQqM3TnUTGbE2CTbh2uQ/+NFf+jhCqLah/EX0FYvN3Dxs5q5Xp051JMty5FdqopQz3qC2TIHBud
mXADyVQZwlCErkPLlpaO6lR7gxhh8G3CCkd0FH6rTVu2W8Hpj3GNBJiilBmRHdt6hAzglxqfnAxH
e7txV9CUwuVvshDXFKnTCcpV5tVsrJIZA1Vhq0Kqg6rkv86JQXsJhob1/iqcUoQd1SvfEvNhzcYQ
OEa5X8IpYNnOf1W/m2lgNxCFGwtERKopTTeWZdZUYYQivsXQZTqbt1/2ZaVbG1FYhrBXiwx5Tsfo
RUhAuceiH7Ang84SV7xvuaUfKsN6MDmxSBCL11mg/62nNXgs4K9yMForQVdkPyxEa6t7Xhj0Z67G
1f+fdQcCTNiLgNaqo4VhpHmsHxgQ5oezXKkrTgzKGQVW72hpJyR2KCcINz3QXcOswpefgNasmuRp
gOEJqFxJcaS/b5qlUoq/39Ve+VWJIPuoNuf45EteK2PlX/p7fxnxyOwkr5bWx2Aqgtm0k0MUduRv
6q1aY9/8uM+1JXCcjiZp8f65qFhpKs+c7oadYNM+ogEt8OaKUXbxVY1mPJdTe9kH4A5+O5p2u1C6
gLqvHucrlYsQW6ujcNiQAwDMXi7GmePZC7gkhdlcAqJPzdMEw66Nhn4k0W5JBrdVgrN5ApiEjaZI
Ib2bMXJKC3fYWbl2U2UPSkv4HS0lurs3PiIRvKZOKaNZ5iPsjS49oYYfkN+oiFl1BKUF2/SIfqDa
K4Lt8v5pQLA8vMDDRKHaUO1U3RDa0v+1UKpAgsr2BqvmPbaBb5Q+tddbWzv94R1O0SFzohT/9TOD
76a0Z0ITOZMFAugyyBCiel1GwNQkEwnMH0x8sLrFlv08FjBdn4uYT6/IZvQL0EZItwxh2H6HSuHf
K9kcaem62O0siciDtxS9DzYVYHisCM0t1PW0JIEBBFnSI9sD18Q4LXVopynetAAKQTOV26/V5VUw
TXt5R+02HI+Exwm41nS2lbC+KJhgdCtEgeXzZWd/ZDyifBYEYzFez3Dv6/N58jxtIH1X1RT+Q+Ru
xDad9rQQ2z8jaoBGz87ztwAhcsl7JrOzFSwfBXVFM3uE7A8IeJTqjaVSMY0v4P2P2zaaNSChWifI
+XwftO/Bc5mbCVUXf2lWvyfIXI59W1I9+1K9vxYzCZRPEDFOiuqbHldjx9/XYtF7LsTAE/BNk0Kj
1E/X6jOCGUrh1FdIwPMEuu/VkuZOi3NQF22mN1GHWC+KykwhI4hROJu6QJsBgNXALPrt4lBubX7T
EmkpkrbxHy4yp6JdNWTbLxfxg2cCIO9G5VPlWkIzKfPgPatBKmYC0YKd5MM+fPdUuDzEoRhgugky
S6aBB7HVDiJ3yNyFDHp2CGW2A3qwB6jKMoS34QxRTzVzFeqj+bbQJrR34HWBh4VZma6JhkFkVg6y
K3nHy1OoSgx7u8TyVj2kqAS52GJDBJDAFaYoa1PPYWVN2EwTsE7RwiNVByZd4T0Pxe1YpfMSTCvO
fKxG6ZT/tODdT5t+KENdqQ86ZmsNbAOsCp+6eOzxQr7EO8aP3kxWKtM+uisFyqe3TeIEgqvnbEyz
brj1KOVDDkW8glTVrtF3MfJb+yQO59IkULH+nO4FFp0iNqWsdOfOhsK7DDzAZwb/vD6tVNHAtYwd
vwUSVzvWy9RRV+iVb7mmoQL4G1X973zUSxqphEBIXVqnGvv6STFSuUsKtLTPdASQDv0MToKV5xL4
cNtHdvuNEAwcmo6CxTkpWHFj/lvAfN3HDcpaDeWD5exy3AE9iUUa41PlVulXL2mJ0yuM2ZLtzyUn
n8hFlXyjrFkTKYZB9qPHmQXWIS0u8Xfif9Wt31LN5xXyAZcbmeltkOXh7jhl24pHEIyeuUNSPi+0
/jZ9yLQR3yqdCZ/AXlCyEZQq5IGyZV/ldXz+7Tv0FDckvQ75TgjP6XvdP1Mr7AZStCyrbPn6/jvz
LTV5YUyBUjT64aj/D5MJJX4fI30FiwoutJxbKTSHXvu+qizUzTjGDdZUYiT1+Oyyd4fU2DcCGwJI
cn0dX6yhK1tFvEH+zhtirorH49vU9fhQuTyICQ7nnuz9VJaKmKjLqz5mwCdlfQe9P9S/HaANiAIq
sDYbu61wi5cmyDoL2PVn0v5cJJPUIEn2yY7wLMfnQSUmatgcU+yRPNjRU4zMFXs85FSH1jp71LE1
kfkYp1b/Va00bcKP890X6vIMn9+hRfB8++gyFDn0JnSZFUUX1i2Y/m1IymOjdISGUPNx6bO66hC5
zG2qNz95sbTPQPxP2nzlvDxAtMWZ+IIbZXiiqQogaYmA/DGiPrGv4XCPMBFUI2hakC+k2auHO0yk
a66XyiTcQgT7NMva7wbE4z2R0pclde1nHzYgzSADPzU9VW4fBFbywMBcFldXJnQ5Z4k93yy3FYMc
AWEcE5M7fhDjCOSfWYYYMu+fSsDmoilf/gnXVE2ZwVQZpwNjLBuNHWTiFOc0+3T6JxQuBLHFLqv5
YNoj8vSRVjtkfELLvNvupjN9QfJ+oBT4deGuCTE3AArrglbOqVVvWRYzj4C8tuLiQH/tDEW+oJSI
vXLVhcaxjidc77+tjspLBFJMmBqRVmQ0LMK4bOWyA9pugVyCAfbSnby+bvlhdApwJzrmDktuYV5I
OAI6K0jjaAzMZm2kUUnmcYOOFKckinlGCVroNSZBqKTrV2rJRMt93gDYgvwEWXbdeLMCo+dFP6NL
TkG3x/5oTRApkLoki/LDrv9xi1OpCHvkFWPCYbcdd6m+RuxWeKchULwP2tarAMS4kYrcOeKQJgYJ
0DrxP8eNqRsOfe1NpfnUEklBiCCCV1AibSlzC4mwN5KkYj1/UHIpXILJXLiwaOojtn/vnu69OxH/
eWvNjfHceP6zcABlpAr8FoWR5pblcrIBRq1vh6iINNX9XJNo662mzoBqw4+IZ0kqEkb6UJCirO7O
MTPVq+MW/ucbFO6Nu+ZzRPEVwz6OYGWhoKKHHN0Zvxn351+IVUlNPaOifcmirnA6n33rlso4quHC
PtkmedjQfaD9ecwklU3pjLGGeFHpW4tKt8vqryOrBvQ0C8GUPI+sWjwTuoJPbTwPmWl2/hAo6NBV
AsokyCPiZ8Jdie2bHfBeIHY3e6yG5aP3aRd8nh7UdmPfbrybGRaos1oV4pDBDPjD3F0gcz1PoVjK
iR9U31cMfu1jXV8ydQ3NXXUylgNla2jpHq+qsp1HZKOhOo17kC0pQrx1Ldw7Hz4RfwMpSaN4+LUD
IjRSCQs3iic7cMN/Mi36NCdrvG8HQq+uXokUFfXzWeovBdIlfuUbeglA57Fi3DWtK/ojYT7SJdYP
1SQw+IKkM6+05tp/0bNQfiNDcL2lu90ulpj80QGeE8Xhe3PFjms4mKVN6ahTvjHSreiSIA4/rTzp
EroCtTrGFCx/1coUNf7jd4hpP7RPVRLOzBXk4yrevLyOxDfiwjx7AZvfg+k7Wc+EUnKtKteH4lN3
aMcVMe9W2v52Jn9G7F19Eyb6S+Wc6cSurYgFBE9hWNzMYtQ46uPvycT8/FukURBSDfRZHribHYaw
1j2zZzvqfj6vAR2jZON5sTzdj01fK7EdBfQRksbb0OMaFyS5Rk1bo2Ut+UjOEe0PZaIKVQfjRPp4
BQqMSTOMFmgencuWOCyLuRXEmGJYk7d9FKzSjT4CfHkjssDuzIJcNDxvJPRdWJW/DvA7T9pwXqGi
Z78U1yLjIgXzyDf3p+ioxrbBbAwTN1ZItt5X7GmYKXao7bYcdeWje33WN+Gs80GikBW7ZCpeF+NT
0FMU2gcP2vgFtwNDmcROoYyxSCNy7/v04ZOn8xlWKTeGjA6fuBUH692wlg2Xk45TQIT1F7yVNV9O
V20eM/5QV+/9ot0aFPgW5AuaRXnppngKziof6lgVYkoF1bMOLTG6DY1/z2Ulnx4b5yc2kVbl5vw2
zw1PwVVBxdlIw4vEYaUIGA1RpxPQcT84btukVZvNLTr3V1t54bW5DiW1mNe1+9TVKKaK1yjk/6R0
IszYSsTkSu8C7nN5+ViU1bY1Nxh1LDrNdPgL6t/SqWabaySrzuZgkAUk88xTrCUUaEls7udVSsS/
MgjASXcHIRag+JTm2bx6ix6VEreWxh19W7D7q1pw8HPGdJ+idj9doXbzI+K8NE8iWIwmndvxECsc
2uUD6hdsgoAL7WzBlqzI/oOySnVyNSyJ74Mcz2govA1kQwZ6dvTlFK8UczKdJxM8kc55gbQBaTuZ
6XHsUqNKYl4l6RKj0pguvkZuelL1ChfuZEpmU/nTrVG37bb0FA7PPf/B3c3Ne7zGAB/nkk3BkBjN
FMBrlfWZEPXTXi1S/lfiU0sGC0gMw6gboNfFdbm2Sr6iSgPrQLdg9y/YuziQXVnAZUxu0QOmouRb
rErmDmdbLaSGUKsbJzidumbsGR+TaI9l1pPAsTgAkEqaubk5I9G+vfiqJoOBhLUHtbCExja4Fo+N
hF5cDr7fjFx/br68z12xLTxOkxQuCtCxvZeUykdX/8Z9oSP2n0pq3IY66Wtx5XWG/LtOObrnsYlX
Fdeyko/yzZO88QzIDA16wmTmJqo3NNpw4SC2ICw5OhF8JDJ3tCZC/7LdpU47iIcdBy5cq9+HzI2O
E/w10nF6PF2CWTvVujmucEVFyXfI2BZNyr7Zg6VxszKlb2iczca50ym7pUPcZS/3pIjTs7LBz5fQ
kOX4g3tNOicdlZqbVcjini+FW0rUy0TDYRVHZmscH8sItfPqyVz4QcQp2hW2c0NToKt4IqTbK2Cz
6vZhNQd60BkVn+67orvXhX2M8k5vqSO6rijb6Fw2AnC9qhij/dqLNHoDQcvLN59ZDTzF8BpDRnBe
03sOepxtaB7ihnIASvIqW3gmoBOCdUEzjzXeEyvrD8Y+8jeJnKMWvEReq9VA+wWw0lSCQdHA9xUG
h+GttY2pkURZyZERs42hiuV5N77JGoWJB2ZhhtRoV2e2DjlS+cDvVqbfjc1qmLGSLv3IasZPI1qQ
9UBdKbSIuX697pzCqPmYQ6TCT4LLMeTe+pXcJaE2hNFwhhyOYZjXlln9lTOKE5cxKJJ11s15pvNo
JOmaRdBKuC/1kwvtcSCkzfU3qOiWTGrphOJiOwAJecVNEUs5O6r0yZSH6MhwtsFTRsR+cl2UlBEC
40o8N7Apstwvqj2LWcLqZpRCsqjVrGvQUypmDoESBLsQnCri32STx+BCiLuhvmejQIIGAW4oKQvF
lHhO3laQOK53npHsNdQQtI5hjcr5G6zAj4Zr+haobS2eh7o6b3Zv8VNPILaY5CJHkLvxJOqyKbDZ
+oNR+9h3dxY/b9L+j8x62VgCPPg3JRvJakHh9vSEStopKAs/wupPdb3dg0weVmPGQMWyEUawZKAC
9DZwuUD2pCWouk9hE21tRf7LM0Rrqqz6oh8NUNe0Clar7Q4uFZR+dP4aYMkb/JDOpz4houZ7kTGN
pDhuQZ2Xo3zuMwKBdW/TrzGBPpVkZv9LYLByIBDDXrytrI1O8uTAABEobNgQrQHc9ijOmtuCmkax
QflhKfXwjssbWHzDBDNk4lUcr0iotmRQ9Z7zJbcaii8C2PldnWKBwkoLvaZJ0Vuh2/KW2NThh6vL
XQVJE3exsWvwNMuAvEFL5nZyJVM0xbsJ0dhMtoY2hCybP+6Zr+BXXqDqPkxQYu1xrgv5sN0k6TxD
v4aPxecIcaXekl2+PCRuGKf5P1/OoAix9TNsb+YIHV+OPtAgLB4LRr0XEzsmJMicSmhuxeSjRZ1x
pvUymlRSQ4fx8u3NBgvpQ4nnGQJ6fM1dHBc4Xl+NTgSosqDzhAFpXdxygZB6RJ4YIpcOuCBY6h2e
iNUjYMI1mF0R0sIEU6Z9dOUz1TnJCXEhbRvDMExGvbGD8jTVuwY2uO0nTg4di5rCG4408toVowiP
MzqxWMoESCO2EEZPpUmnx3q3+7sPky6fVRZbmFXK/B0mhbp+59XUgbyCtXBsOSeTfKXKM/JHsqhU
s5llhMkgD9tVCDgNEdxP35r+RWAvkRVh1Der2A/bKyiCXBHsAYlSToCZV2bw5FjDxQaQ9fLt2kLK
vdPJoxdVYlvyV8KWALGFYJ2NaWKo9XkZA/gQCOTKEGdWEOjyRoNoHnTXJs4hQIW51qAA1XT4XpBO
dEhN7I2v3O8LgD0kyDHiwTrfF/f8o/LZ6tw7NbUfe7R1ZW6OQ9NQz6uNshHPu9HAne6nVeyghKdZ
n/XjvVNxvi/SphTOZVQTYUcziNoD2Xw4bTcgS6mNmiutU2GT1JQCRnkXe9myrvaTkpsQvULoU02c
RQukHErjEgVh+6Kn3owSQVq3MVuMGcvCMAduoTyxmXhptkdycp1aKQUEgiFgCTSMN7PHPXlLcVk8
jowDIm1d0+JG+HYt2GXtEWV06Pnvr6WzAJQb3n4EL8HiZq0n+ItHmi2oT+r1oCd3lRr9TVLfE5+n
zTvsTW3a52JVt6F8lpcvHB2ZpbIg02hXhOIwQW3VgtLYDIk8HGIYvlJXs37dmTSRnMY+0ukeg0lx
6kAlR87oeH8brvcJn5FWTF5jmv+6Kab29RHe9sdrMSHTR/SlVhyB93PA0a0sNPkmcndmTbVT2EoK
rWsdCUDbLWYtNY3ucLMMNht18atDwjeU5Gm0Wy8WUfHiMm3arOXI6mQupRc0Vwd9kZmiSaIyAvqw
sIN5h69CBAtAtWHlB/de0WMumoFs68rtEY3xHYZ0tiZ+cZhJ0qgSdf02ohw1uOf8VcqJ06/gO30L
XIixua6LTpO82dVPxED/Hl1L5DqyHt+Kg617lzdMVTxPaWPcu4Q9y/6QPXrs9Vjy/aaK9jUWBPE2
NYiYxEfa27I+s3eP1tqv4gsSdIMy2Ac69E5CIeSZ2MHiC3PXS7ejY/X02QxgvKFgtuf8cv/XIZj3
vPrt+xoQ1UpEoNWYADf1+qjBk78DwtqfG4ozPmjvuNUSm8hhTZX4Bfhm0qbulB089evknejGI4lc
YhHQ9WB1hbJDLFamphEc479JbKT2c4htDSFNPfWiPpt8O0AHN76EIbYiDfACLbCbXMxSIcsd+rBG
dajRY5Ddeh1Bp0IFxExp++2D3rThnVK1w+X8sRKPv9iux3i1PT0q0Ff0xN5V1EiIqdAarzVijHh1
j6qslxAu3yUfZ6jiOGLHMSrZ1vAEzJrwOPNGBA2fklhil1c0P4zFVdfj1N41IgHvXi+p4HI2RtbA
iOixrB7ghV23b6YrQFFUyDGNYcqWK0mui8QE96gt6UPyIRXmp06cgRTzeXsTUXPdo88WOY2eLIFq
1RE4uKKvssPbiryvXvV5mQZmKYD/o4tnAXLxRSDx/raBP8kOiYk/uQs5bAZBLtGz5bPXTgsqdEZV
ATETc9ZkuF0qbh+VyC7aj6FPEF0OwXzmcOOOeiMheEyLy4IOTUyL1xRZzV2dDweaT6KcislAXBRz
MMaZ9VM7/0gg42719UHdbsUTqnNd5UJ29ZMIQu+jSGQbCUt7qQ03o560KgU4TzRGXy+mv7axl8SI
2Wfo57Z3cYdlycQLTCj8rvTHvg4wT4tYoMZ8UmTCyiA+RRIuRqotAqfrlxku6Sl6CZbYK4Gzuj6W
LkyFILbXOvmBIMECckHSeDgZbQHtPgWkZMIy5NPRCLQkN2bngwH3FKQfVuUph6851iA9UQDIF400
zm7Suq6F5J3lRra4sHK8Wox8PdVfqbDCq8XyidNQnR5qFI2aWlgdooMm6EfdlZyljzplr6ZMjoEM
CPIgrOC4eSLo7OPWxQ3GlgYo/gd7MpGHhJfx3oAUiUUzj+kQmgrJMNjuzzm7kx5qIT2qj5vlmNdT
3CPNwrq0CuqalQomNAjUCB3ESzhH6wZ7fA2FrTagnBWccLj5UzdsnHlggKy39XsPdDz+wy4bDVdY
uG/iANb7mO2h1nvGrhzVC8J61epOc4PFbQ5AYmFVbLljVdQlz0uZMskTpvTsbsHzi+OKImrnBt9J
o4zAFrKRcub6QAxXgpE4uHX4VoIoyfk4hVAyMQHWVhSmKRnV5Xq77/SS84wW16UlNziS3IODSMla
SEL+7WTmI3a3mwb9aJPIwErOgk5j1sRQDr5VcBMbGVO8VwJP3CXycL1uUEesAv54cvBntDPBJyjA
ys7FJqBOSqgJGTEMdHF4JQl5D0qPHokkWKMA2kXYQ/Z6tOg5U0NwHtKjYSr3djt6gAJyHkzzmVUP
LWz/hLZ3jNJy+G23OeIE13VmcbVN229t/UNvn7aIF+mrt+dITlw7svEsbgyeJsHHoyq618STKYBe
xSYa4+OAHGJ9S+TGrDpbVJ7vI6TCnR7Hz//YQZ/W8F3OzlqvWFD2OLela+BnGSd63bPEqdc/tbE0
jKo6K6kgQoQFvnUbHdq2uAHIpisy6hNOaGpLd2tGF3Ge5VZt+8At4cJbU1bpNs1vBYFSAeBMnrKs
9dyBeIkne/V/MICgY1egvNQK243hgUocFigeIhtBblVNcwZrlmxrgy//9O1yAkregV0FHUCTueRq
WBaemWmaV5ydr4wRYo2jDlRatggr0JQClDPLfbgP4C3c5d5+moUhD+XVMfxyDL2Free0PvZHEn0k
3WhqQqlUzk+QztWFL8JeMGFhR1kxxWZbpU7fByLSR/7wG0U2hqRIJRElcgl/u7vZi7X4eG0AcTeX
SfLbSdk1Mo3zN9CElQEKS5SadXWRE+hZyg83YQX9aZS+xFYivZsgJp/nTGfvGCXWqxaQdW7wuLFS
c8VK3t4oTmpA3XZ3ResXACoeYf+SiEuOgcumbBzSTsSAPoLcuMBc3jQVEVoR8IikOTspbWzYsGQ7
vh/8rymTgzqn+TupoNWMkVrYnX2lbCED7t6k9uNvegU74KXvuIHjRhb4kyeZPPabOz03UEE1ToX9
XCLMmkG2Iw8nZN5P698hlgfdct5viQLxfMF1n+MTyptgV0PjfEDwh54/4f4mSpOXkrhGjDedUDI9
AcOBcwelHSK4+/j/lISisVDtDmfHO/14eNAx86eoaFqs28riQqEL27ddpxmWrBvfpTWHKjnP+I59
6NFUPF29vnpLryIBI5FVCufK4wFQaAE1YE9iH4Q9Sd6fKFXJTTUKGBgRLnN1LTSDrCEkKyMXxqAs
zWm+YHDlxMwEp5gUCgR1j0P1YXR/MhxgSjxWL+m2rQ5CWBbb6p8Y1jEgVuJWLMkU5UHKC/ivvKTQ
2EWpN/amsyRbYi8p8xCCozE/1CNweZ13z1tc66GVv7yqAcNmyJJJzleTa97krU/v6rGlhAZBnQBr
I3l2ZNNU53elQJiIp+N4b5ZZgGFaPKXmXL9S2zozpH/H4kM1QBW2heViiBw6AF3o4bsbggRs+JFi
mSmQfL/ARF/RH2R09M1mRyfH3q47fQ0GJwRinOAfHBLA/hH9Pgqc62a3O08ye3srt94wavbNFhDT
O3MpSDoXeMK52pXkZ0H+GZ/brB03S6NTFLJcapOWCYTKgSzeHejdJZay3qvuQPT6LVIUjJd6wFtm
bEAqPA5nwDR4UqDGcjG5BnNXy9nGVjNjsDHLc4NWGm5hqEDCXObQLLq5tUYTKKSpH1rnc5dAIcDT
Xd9Mk4aqZ6OKP15eVgBLcVlOywVhmOvboxni2aGPLPH6+JTxeRBvpiaz5McRurfCl+VygVEkgKYl
tm6ELncWG5ZBcbnDm06zPo5J80Z+1MFyCGPgEjpD/y1L9Jx1WZpTl3zA32rrQN+PwJG/vn94RlX1
zupsCo7C+prpHqmaXDqJ3jmy12tmXhfpuVoMMscZm/Va4RRXpOeGuqjFhwdr5sUitFskhD3AbKCj
z1Mc1fArbhKMPHVBpv86FxSiWPcA1nSk6ZbS+IhgpnHhH2bVaZrv2RfHgBy3p0s66zr+kWvzNNt3
1NjxzLQHEXUtfMVnwLDYPK17uQq7XQBF/Aq2Sjcx8To8pgFE/Hi5RsOt7yrBnTo7oxqefNqfM7dU
4YpQ1B35Klz1QQjljd8rPnjag2Pp06FdY1x0wohXusNvVkT+9KxFMzCKA5iFwE/oQHhvWZKcmB7B
QoA2K2pedIHSI0hNNGhWmO8zma8Xz2+D7QYQ0fWbBSKNjl5pq2xUH7/ZMP4HpALeXe74kf3jAJM6
08Sd+i082QCtXBhfHcJH9gf1TiigbW1INM3LCznDhPO6K2WzIWpFVA32jAdtJePsBSFX4e1vtTD+
K9OuPHJ9kp3N3bO2ScA90UdNFrwNLLjHtt3Twjsqm/q2uvK2DjzhR+FBLBx8RqxSSCXpjH9rj2yA
09nLPJI8ph6QcXolMWTjFxTY1n4cUeTBzE4I81F3qKuk0hB6Hnayi0cXwjGyUP+EY6MixnHkGeno
JwagBOoTO+Cu/AURuaG8dz0ZiVsXFo8GdiYqmBlzraxhs00Zy6SJ9K5dauiRcM+QMctFDqfpN3Yr
ILwv89ZdZJHwm9I+kDUri1AAMHGL4UuHVdIEVJxnI8DeCVICpjxbygof2X58bPya+exUz+DlpYyt
iiYelhIVi96sH06a+otht3ZpHXkbHu5/O4uNChqz6Nb9mvvyjLEAua2X6zbAbmtteGwFWCSnEl35
5yihNB2E5KKks2mk6qXzddR4c7YLnc8465gP6fA+ZSn2aJOAEkeTwCFFHcp7WDb8o57NKWb95ysq
outfNFPF6GwIKK4xgIOsrrAFFv/D4MxDrbUfw8MIY/kCmnfTjni9zEZSOaUK+pm43ZJmDCahMnzV
+ph/DCOAYfrxwdbMZ4w0wbpGWvtTWHmR5Y6V5qmJ0gTxYP1qQsrPvIcrEjwxYmA+7q/TD0EJsGLi
tX2kXC5/At30kLEs/DJYuKfuxE8Eq7ipCO+vFGgjcQy/UxBsE5R7BHGGO6MBsrw2UQrOvSzYRHhp
MH6sg+LFvSTh4c/3iGeUE2oFe7908SLe6CDJmLeViguiL7RLTGuxcy3mgpx/VePLcvF3e2+rVdmf
cnDBNwV3ba27g+cJ7p34i5wM3g3UThTr6vJP3nEU9E6FIeKdG3sx7vOzqQ3SRW4gikn5cbnzlqMt
VlXqcYODK53BHH2b6uETPgepHW03v8Dvzmk6c4i40c0IsAnxgvJdzPmceSkqCTxqhQAaC57tHrde
/Umk1iSXDREgdc276gdc2675+Mr/0nUPrwtnFVNmm+bkUd0Wp5aldGBDX9DgzUiSNS9/5vDvMuRe
RE+Tcss4N4NRqexiMRqk4v9/0BETgJBcvJAX6NujbqRgCx+eMFaT2bijaIy5m3NDap5i/SoZvDQM
Q8dlnhWZEJtYCkE9fOkNpwe3eULZO3nF7XqPvAFL0yMh/2aqONkR7O5I6GHOaRSEsa4fFXxQNdTj
KVXdckr3M18jCYXtR7QWxAT9rpLlgDbSFWK+UedPR2CQH8gbE3NBTCeM+uNCOYb/gBIAjqKa2R6l
Ayq8H7uKDHGyiQWtX/GAolTtLyvdF4YSRLVi6ZdW4WotcS4LqdayByakdDO/wPUoZe1S+WKpqYeH
23vIGW7gWvZIQyN3IRt+e7os+vvD724bR9UBr4vgeRKNQJtU9DAqk7RLxEDx7Z7cLydUNGjyEPOR
NVgs3SY6SbzYBz//H4zoT0iXsv1xr8jHlDFk9LUyuCXAOpD09VU95RgD4A45qXoM4hJbBrZyHQu/
3EMOMECZcvciLiNUw4/GZagqJh5D0zM+LpEHsh2JxuZHniHInf23vn7cnR5lMiMb5RpgvRrMKRHy
acHYMT6E8SXpB2cDDaidsHte7rRWmywp+SU0g6TlRRgNj3/5DAp05Q1E5BSqUglqnNDouiHmjJz5
Ea37cGVErq7pO21b+bStyIWjfJsG/QtNre1fQcK+HRXgWdfYuDHTKRkBy+lwF7EarEQ/WaauCDbr
k6W9wI2f9TFJmMk8jLPGZIZzK6esuaGYNK+u7Y4+/hOFbpfXXVyl9T1YBxEyHDmTHuVfwa5s/ogH
PnM5DViJVQB73wyPgueXM14qDYJ0wMA0NLA0IlXXL/RLt7esRoq7jjyjHknm+U3Dt5s311tPPrlU
u6vK//Cge3IXQfqpfYuOpr3rkUI05j+MunqP0pA/5hNonPZh3DXasoh3RUipSTsrifyzHQx5bfyo
Dc1moFrFmyQsHZyejhwuzqM7HAVluw7NfYTOTrd3xYyDIN1Vp89TXGHrkOD2p3BZx+JmVWvM7seo
Y2yqDR1iw+GlnzwmgDCy/La9X2oBgWD0DwonfNtfWPUdtxxW8Im1OUggvDEtn8Of4fgWUqDkJC//
A+OO2KmQNZ6EpAGRmMNjaedlguDnM7VXKwwBtRTdKOFeKANthkiPPSs/rHgq7ADzrhdZDCB+mRGH
a9H9hfay6eiCVCpY9AqmeGpBBUpqTYHijz4Ip+dAh9uARNGUBx5eOq8wWGLWc5a/v3FlUQKdOnUY
DT39a1Pz4X73Czu4yTbGCde1bF0DOezFZ6P7/wtMgr4V3U8XGAGUaBh12oFN7oYDbvh1R5JxmMYy
YazfvxcMaARzRWDruGiCtfryuCms/4+lu/XHTgNedmZP6mIk6U8h/kskasJOWb+SMuU64YybW8H1
0Qw7kgi4/OQXlHiisHDE4YZe0qc9RPr8uoRMK5/6H29glHKI92VxXC2JQkTgsZd4xYFpBDx40lcM
wlVFXMKh3/eQyn9o0dGomnKwhbhCIqe9Wpjsl0whEVem2k7ccziJEtbaLt2b37H//lZKmeuBkDuH
00eIjcC/ZYIZEgy3LoDzW4ldCYOK2eGn23hr4uZ/A5QYZ/ZYk8q3v8UvRn/uy/ujjY1E3aSdrSBa
jw78Z9/tgbEwOtF0DCJ/NVoJ6G2KiahENzH5SSQgVTOvZ1poGsuRMDps+0eRhmE4hFtom0AiE4BZ
dhWTQ0Fr6v6mKOfWFx5TDZwD1pb3PyNA0IipIVCvRXJMdOMxIRJKUKCQ6fgdl2WQzlcRkUKtlKtz
rUe4dvc+WlVYFYX7Ymka7SyAADw85ElfUEjBXIak285dtn5bo/S358wGaovXhexEh+hi7yeetDqL
WJXclVnUSXKUEj4U/pvAmL4dK+92/xkaH2xVhtOglb2why1W+7MGeABjIy94amJ7YY9SJlLl3ppo
AMRlR1qHNWcIdgIjH5RuGg8wDsIcnSa6gdta1qbMWUxtlYRIReO+9Lc+njzSXVxBkD6a4+eN+ZGi
ELdK9b/4tKAyQd/LT9nGNnSZG25ai2Zel/DG3C3/MdgxrRByItkDnMSHJltNp9mI0FE4Mb77SuIN
DFwPr2RfjU5we4jsysTAp/vP/wLgFJm937ueYkJA779u0hFqUro1XDlxjWexHlH6p0NrwYmmNnz1
Fq1abcsaLP3N5qNUF54EhF0L7akrsrngqRQnCmafp/D2fINh6QqTESUQlFZ9hdwObDkp3nB9JZBT
mIr9eLoiEjMxKIUoRJcl9IT/BvQTXy3qQVq1UK/0Voi87hx/Z+LppoQYS76/o7pIuW74vC9hV4Ac
bKhihqSQYabrBlpyL5q6ra/LU0tHiMH26E3usAzsc4rXboqbtS2jJLkBmXsBZm1rOoC2UnTJcTIq
QviD/AiU5MiULeud7HCLyX8+lpUQOEHTwe/PWhEZObMkIXaLi5D7T2IYX+psfQzxmvLn2IEoGqQ0
KEpA9vwT5fqzGfsok5PspUBnRxBHMqDzwYXlHWbfN/p5tIXHQOfCo1dzxujpXcbS5f94gJdmIxKe
EtgMBYiLI/Xe3u/ul2tjOtF5xM5D9OGRPcgqR2cnQwSiqo+obAXfmFFScRWTqCHs9BsQ2mOO8pQl
iMOBe66L1wJx8A29bJBVGY4caITVcnR9AxR9ceR5KabmU34CrrE3TyHk9O1UC0AEfMUjFxidlK7J
dMzUv/YYaE1XiOWZIV2dLLCgM4csrKc/n1hVF802d+mzqkT8fYdqu0mTW0/BHG7iMdxl3jl2pBJA
Ki7xnMwviyTUNbLUQqnCWGdP9+ZTmdBhalKlP67dLulAssCfn58+mSWsoeA15LOWwOv1YMrhzC1t
3B9mj/fPtW6YQys+by1d1Vvrs7YShZn7UMZPuhRuKAo0kSBTkZjScUWvwzb5f9O9vyiczJEuJ5J2
yQRSdvRcEmve5kUqfWKQDd1aAubzpKaZhTaCtnRLqalloa/F8a88GjSx1mZIwFbZ1QYcz38N9q5v
L7st+/v4wu5U7gcxsUWRF9xX0rh4ydQ4FJ2J3YEKfn5jTMLhlC72+MHRvuPgbmMMt2uDEajZbUUi
IAhoSgP5Osu6AZN6g5SMUdS4RnKrFWUeakwYPx69M+69G9iDOosTKHSqRm6f73tK/d4J4uJQI7ps
LgGe5r/mDopNVpO83JnykaZPcSWlJJZodV+boRNUWjOcGvoK7b0+Q1QPnw6WKSWCGEtjNbZ4YnIB
tmXAsNuwf4e2hr/q0kgaFGl39/ru1Fpayebfc/3VvAxWro3/JDbOhjVj6lT0IE5pvmdspRZCP8Vi
Nzb1+fzAQ/b6eQS9bmYpEfTjc+oIoEx9g9YmIe+ITRjbe4DPoTkJY3nQq+zO27XwdODmS+m2TI/Z
vhdc6gaCRxfN25PgjWDFvpvqD+Yozt2zrZTQSWeC5pqBu/h+arxliQ4ojp1ASP84TnIoauM9zAwA
vjjn8XUjsoMRIrG9UJPpTIEf1Hu58DVZqxG8UNtkuxEK5InVxwH3iPtDopMQys1aIEpcEqHTyY/e
+BHfI2Evyua/9DNDXZpVUjr5qOJjit8lKhTRoo9cdP6H/K+zURrJVavATdkrE8vfhQhnFHNEI1Pr
14Luc18tARg8M95GznUIg0h8GbqEKsZiJpoQa7yO7TjSPpnN9KyzfmTfG6qCLP+9wpnhD9lYW0Zz
yu9K75NzrPiHkZthcovQnsTcqsqGcSkGFR9/wRVkw7t0iKuwjYtf8hKsxzAVK3SZdSGhjGdwiLSe
qtdxA5D8pSrcdGViYJ87PeTKFPF2ReWE+b6D/95VeyWt04nQRodE30s5Ywue26nWdVzj/+z4lXoZ
Z3PzD6vt8PUlZvjAejb/YXWws/HOwAe+pQfXE/JfAyLKeM5YI645ixHye841Jsd8DtMiqjtHKVgi
/x5u1g1bK/JiKi4ObGoduS6ye/5lQW8nmT+9H1M4V2SVrk4ViTICBoxhFqZE6nwbJVYxWDGKwG0Y
0XeJSx5gDG13RgrUw5WL3/Pm9ixgycJG7p3uVbRsr3nJhma+7oHUzOeGpdsgiu5l5EJCLeQDVOtZ
G0SmU02G7ef2UtxtYGpt7M/Mmc/7FPy+nT3ihszLiiikScaTAbE7b7y08v+PjnuxXGEWmZmPLJYc
8X/lZ0SJUj8+px9pmGoDDppPOMyOYC/obP/tGgCVXxvlTWiZ1x8VZuvhhaHrhjY8INlK+YS8FjgH
R0S0aUMDdpOvAUZLGlzlozJ4eQQ2Jebed6yKl8rmg4aTKa2AMwl6cC1Zw+/WvTz1tY2/T51T/DxF
Q/RxX9swD25A6RdqI2ZnGT3xOeZIOdfWy6p+hl376lgD8JgrZTbau45DDsGEgeW9DKYMZzMbPSjk
70BETbudMvb4VmXZXbd/dAwnQV2qZpSSLZkbCJfTfnLfN3/m4YGv28TQXr05AqHLwkP2UlsSk3kC
U/OtsXvWFQpX29C5iPaRCvCcBO8IEaEr95X9lGmMLhNM69vHIsqbbtyZUl0nBfPdxk0dfR5E/Mil
UiZdrGodBPRgYPA7oQ+FIBYyXJS/nzoD7zhS6GVsvOcD22c1hLy3cq3hJ5T2jc1exmnin3MGlkn6
y4nKs3n2KYmxbd1fBow2XZ4nZ33sdcxReRvoftQYtnGCRZ+yx2PnYuWW2uq4UzOo/Yu+p6mwQFCd
o0mrrZ/r9YlmtUxaFhMEegmK+cadzOqvDZygmg8awC1LdcUiBtYZXryAweW2Epzy+ZZdFIVFe+1c
xEaf1H2YN1OkTMG6ddfDWEI1RS7cZIMLFOf699OltwhxV1MaifQBcGagRFvonyCPfXRj3/XB7YSi
kURFoZtnKvfXtr6pJvzPk3VuFKkPuuDETZ0dMIXlnHJqYXKtdvL1whqvzC1pVRFyTjONrPP+CKEN
q6CZmg7APo9kdO+WEo5OzGF9fGnVO0DH7+TLLXtFoXJ6GuBnRJh6YfM1bM5vYBzyZh0CbVO0nG8c
5vuN5vCyA6H8R0jeQFkEC+cCxWe5n95r9giQb+HKqh61lrnf6cBx3UmP0uigf6uW9ejoXyfRuPI9
7R170c1O1CbXvcjbma1+1UhFn1TtUCw1CO0ehIicy/8wJ0vAjT+tESKedWr5AyHUWCdfYSEgXhhA
CUsc5wMVy6l3RnxvFu3EGyR9/dz3lIYZxAThswdsa2pjDtEUnPOzC6/b9ARETLm0PXIE2HKTFLJr
gKfSKL2Vfjxo/q68vQ6Yamzp9yS/+hrgWy+8AeWAfS/z/1FJdDySKAIPWAVlPeIkZu8+9faXkymR
tBUSJs4GSCowNdABN9zXENP/1n7oB/s8Sm/cG6B4UoT2jYurS8OzsH96/N+uAjpkfgeVaGmbpUF1
kjg6hGwB6chUET6m/uqMau1BMQiZOxjgxO5t/xZVKOMJu2VI7AJQFBpTTPBgxIzJfOI7bR1XXNEj
Q/W7YYxQZzczoNnpX0i5hr9OSqmo8FWevoOXdA7N3wAvCZ0jQgNU21aL9eCytNWK0vNLccR6dNBN
7HystXHL/biSxtqkcFJ+aYeEwohnMNgLza+sZvDNtjI2nCHLY6JERrQloZ992mPJuw23k8aInihG
Fsw/2NC8G7okTdbt1liyaZFKtvBOAIgMXVTPhOWia+eVY4INYDoYxuvHETJAarHnJAHQIs3xHZ3d
7gY7QAKdAEDvt5ZxPGPVpahcoa96f5sKdXw8uHOy8Eb0rk34JEEUBo8EAEt7x0zAm5ySSwO0jpat
zn9SFtSWzi7rO2OWajtKxn5JYhvjrhIxlqv1dHIOccmYcb0OEWu9V+VLJ+Y/pNLKTQhyLbikH7cb
c6rFm2CnweJaQj5Hqa+4fxigOv8Y8lALavaQbjYZ8HXl5ja0FGjG+4DDDrl2yk1YUCpkPYtXCBqh
7lPcBlpbags9i8dR8ddRVRLMBCXLcjSRQVn9HwRu8EpHMO/iXf5OqouR25dIb69Yb1zu4fSAaVkd
GjRvphubnH0ViRzgJxtRMJHkHirFIel9y4Ih5dbzuw7mrwSgArC9vK0J7cdNhrkegbscUCKrbqtg
UjrhKCY6y28r2zk3pO/thE6CQiKjPkc2S3ZvhrM3uLl17+hba5c3SmDWqjShGgwLJnwgbUYiQrsd
cVvC3TseeL65eUub9V26JNa+Opq9zzZMIDDDJm27rQxC6KKGxA5lwPvSJ01nxWZTr6wYZ81tom4S
M8VIsQZNRvlKs+f3FTHUM10NVvozx+0Iz9WVoWqxyUfhRf0DaJ1yFfBBLm8DarVmBT60l/zHmBAy
kpIl+bKKNkUPEQPkSE1StE4wRQp3Q0xj3EN5SW0Dj5hL/IyFHXNvq9amwM2kvcxO0Zok2kbQJovt
+BfvulYn8xGQ+5WBJ/pLwPcwqwwj0aYXFOkpQMcP8+kSFz7CYHVQG8a2fww1k4mm8D8gNgaMlzxl
YQEj6MMZ5/GYVvnQkyNyx7W0mA/dkMg6gMIfcfUtvxBtjZQK4tiil+eYbnpD10kAWeYRERcl8oAW
XgWuoXwBrnJ9fajpQUihMKMNHSJmk0jMZAdmQjNDYhR1HgG+RJoWRvwNqFlA9UWcQHaDlfbSJZj+
J2/lzwTtQ+cZ3Bb2xn+rBNp5rd/HWLlm7O3wrnILry0S++/4ENy44ZXUz2b4nRzDbtwLtCO8M+fu
oDXzs97whneePnUfSOjS6xsGHhMF18cofMOJdnz57Ijh8CCNBRzSXBmPWyGFWAyFlWTd5/nOrGKe
Z6AZesDXEaSYA9onK3bGw+TaW5BKkk8IH4XtYuOQHfmztJZMiCYQ0CeFjbhPXjWpiD551ehVPsSu
KAhdpzZInZPtzKkuscij/0VkHHjBDG1f9Hpz9f+9GSeTwbXOFsYouNUTWFD4Zl5DRyn5bMgNdQ3u
ePFlLZFACtHiixatnaaExD71MC57F5e+4AWisfcwUWQR86lH+3ZFlmAEdxGISdWh2U9rl0RsJJTt
RyktKgZvEYwqibwGzABTbrQieuJHuYchfZDr1nAKwGMw9b4dn8u8oz5D3xhtW2QA/zuip/ATX7dB
6irJNqCIEejd+6jcKqM1h7/Y465lisQsHVtypJMwl+ZFIn+Q2vaua1dZOM4GMCypnUxrT2zmGasV
Z7UlOueFdQQxuO1pkNX39wRYX/N7PzlCWe/9FLi19HKyNAU482U0FsXki2xjcGgcMu/OfXI7gTkz
vtBgBmXTo5NJRp5AAeXi7+/zS08TtFgV174bnJEskBuOdNqSvfy7mrGnDs4wozIjDIPNKwR0OFG5
XVhMTfcNs8nh2V/SiJyIH17zuSnXVPE9RVGRHVHQ8VPAaQEIsCIw3RPAeC2bMfIVtgzyYfHsk9Ad
NSkC4fvqKYpYGaWrGx2Hj7J9z/124WErcl7HK6jk9WrIKG0vcRWaeGDH4/qcafGbZwE2C98f2Sir
joaGclXPYcOeYVCInTD1sxL297LAuP/9ph+lpBcRNRnbmUHYk6mhw2NKqAsEzbn0TWYWhnaoQ0Jx
VtX4EO0yWXRIUJgWWyoaBwLnDtuCuEdmysUKk19/IiUREJ1KDl539KCwUSk+wzYuDrX6GD0f9NT9
PMga4hbNJWC7u/o4GNhH9Ey4UMdQ/Gup52dxaZb0eMp8mAYHeHV/sI5wuw63eZz22qv3UoiAxhWD
thwsp4STnntz8kLimp05Cmn50d4oyxbFB6MOme2CUQHc1gM1L4Ef7bukveI4r8grScUrZO5+KmC8
nzribvCOoNzgHg7FTICnldUTlmmRqq2o6mub91bT9ZxU9RGpNGchusc9JnbqDbFpw/H/8DaDuIFO
jGYrihIxDXV/zHLQ2Z/88e0LosrL34DsPFjesk8HAoYba42QViGtOsimCW98HFu2RWNlZXuzN+mS
90KjHW+OTlWS9xCwH+Srzk2+e8u2pFE/uFNBAcasd8Z12l2IHzTIpdGyGZ+B9bdAK3Wbz2NK7h6q
+XSsVm9xcDNaBYQk/PiDF6rl81fgJ1p+YXvjGe6Hn1gvDwg1FZ0T/WffcqBHluaJVhuEQZbIlv2I
LifpMOXt01kUkzOf2ZzEBvkkNIwVJmTvKVN7lUEOMiiFt3GCROQ5xiaW5kyZ48Vmx2wzRuaKrft9
wa/pwcEJJpmPT8qZClFsc8K82ZtQ8wv+Md0eNu+cH9IZQtrAnAXsQ4lStKro3eQcerV7ShpQIeHy
YAUERwF7REKB8c0JIHCErFCKn2kcTwezihkxEL0471tMz/kbTl4g+dKrac5qC3Q9io2kH3OUXGAS
hRRsiBwaeLhhEv6Rneu8P3qoBTY9xQ8ipbTi6Msx/JDsqYSg912difrQJINab5bS3yKscaonwBMS
ldE8c0scQm+Z6XQgm/u5sSEXDJPMStLtRm36CdfkXws5mXMMFCoJE7FdO02n2gBRl6zzcxcWW2A8
zyF4aZJwBHRPerv/z5bmtQvmqf85TzB+i8dE3hhACicY12erR7xhg0YFl2Qf2pR43CUQcF3Voth1
yz2trNSW580Ao6/V51QBHvq/yHlVARJ1oaRmubp2dUgiFJ6qgcfPWnJvz8yfzE+qnbnyNT6Hwz07
yDiFfkzFLnIrZljkSUqiP3eu9lBS6pUrsI42h9ApMAGTlbuhVtPJ7HUdRlKi29dElxLr5YlXOsl+
YIP9jy+C1ThCM6YGbAfc02fnVFpM7EX9Ga9jBcl619/qQCw7WSnLQezRa2DkX6/UbKDt+c06yrhL
SU2M88ezZaR6fHk9WetlM4Fdz3BpYhFwAceWlPKhDWZCIdMs/xdOBhx17LAUjem7mDkQPgSa+U2n
yT/NXQor1Wh81+NecVMrnX+zSNS9jECEkCgJG1e4ZPCR4iUPW+z+BB4/Mf6w5liKMJnhSXm9xvNO
VCM73EW2FgeO0NsYRA+qdxZxMbt4RH3UZcHTDcf+X3kT3LVxJguSwVzios1oSLamysTyyn5d9K4h
3KNr29neHsp7clVvWjrYxP7MSdmO6nrmHnzv2imUfV9FKr13lrxpUWpggksfKbpY6lpqHcZ0rpeO
L4ld4TvyW1xK5Twj5S28DzX93taeBbYKVTdr5mcxPyUlm2lPxWHyZXPTgmaskaHrWUPnRd4ALduA
1tqHiDRP2KFJaM8Lk4odMu6272UHGWb0pC2sbMq/lz/cNPFcmNm2K2wM2gay1jVkhf/9ikSvuvwa
3kz9nX1IZEpobmLMk5+Vi8GpXxTMQmaMzx6gI6cSJR+moOldyJofpAhKgD9vOJsD/I5cfJSFxOSF
eBasYFd8ZX/tq279hnAxI9Z1ZApgF4hTNqHAn3SYUdUe8dK4lWKpipbqj26fihOUHZmJjHWSlGkY
X5Gn+r84f0p0ZsSu70FPW/vrOMCmKkU2o+MkjqAlSQONLIdOA/iwiITD8YvydTwYy7t2lDkPnMIc
0bbxF4fBkb98JPUueBgZdMjGQ8pXcUwzsJDrECVTMGVNfss3Dd6ztJo+PPPvF0WkDpq8e98IYoM5
iYy/QFeJak0Mqtq69Ksq5gmanJ31ez+W6WdMjWtUsr4t05yecona/6OlNdaDbVPRtUqfIY+tFFK1
wy/EYyDZ15O8lFaBfLFEh4cDDv71i6Sgn2V72brQbAD8TQsgrL8gyREOj7exa9qWNmwVe3u00ZXX
A/YHVO4Yv2rFVUuGRHFNdOeutfx/9kuk9Bnq+nXrr542BSIR34T4vWs2bD0mYiProf7/jEs8c582
Q/H1R+5/4zKLY6Uy853IFptcm4EnfDdDB71nj6WC4T/bw0e10em9ZPhMWH+Un5rf+LN1bcC2PTPl
XrDZHgqhaNmBy3U9Q8SqICahFKs2bM8T1p9Gecl2e5BY0evPxFI/HPvPqtMs5uIZ46ux7o4FDntr
BdJhvQjVVb6MuOpkeOLbd58AHcHDx/NIUMAcSKi9KgsrC90/qM6+d0pcDQNMVAGbYwl2BthaG8Wr
qzUTaiL58P4NSORUHul56DOG3LlVNM96ELlDOQytjFGeXq6xgOSR3ny4byrmsNm8n0QDpzBvNxRM
dvsqB8EYdH77Pks3Zvx4iVfQiAQxCih0Fu4PYQzhgoZPX5n3nlE+hChenoe5WATfztIekOZoH612
DKIcce1Hue4tZg2Zd6C8glXX8xkMvuTIGn51TtPBpJjk0SfC6gYzIjnD5Synb3Dhz88H5OOrzB00
vnRZBhYOiA4svCzI3SpYJ2IkCst4qExSSxsQmCRk+w9jcKWoH0JuGu5yfIE2CR4VrjeNbSsfVG1u
XVE08MH4YeyBV/GeF5nMkF0wZkMwrqcoIGIsXMFN4ypuAjkqYblDSKNtIi5p0gNZ84h9etMjorRB
uQqOPZqL4s2JDqQoBt3UX9d8gs27AuNkUMgSRTsEaEJKN/VW+AO8Xt306WodsTwnSagi+H10SaKi
Kou4MuDizKx5NXcPZblGIz77Dhz3W4FSWclEFWAhDHVWxzRg65z23a24woiXHNHTDYvyuQTo75T0
Xsd0U1lbwg/DffcvxO/AhPWzoTFcyAWNpUtaYim/4V9z63fDx5vN+I08vWx3se6yJp23rkuNEAoy
vh006+w+m7EJFaSyzC3XH+KgQknS9KTKKWI71H78zNo8+b31o1TvU2Wn5/tjPFs9iArgjhE5wYii
OyAvO+1y7rxRODNVySMcZkmMRoGuqqMLWveBS8+VJW2hK0+wR71PGPrP2iTehWjV6dciNJvayyEO
subIZ24KxB5BSwLG1YdGOZ4xmvJSjN+xA+qOsVZ/Y8oY7t8EA26Ol188cFrs+uHqEpFnYqkXuv56
xNPBIXwJ9N5ODFje05JJRIYnkWbfGyRXtNjwfY7xs4e/Qp30PpV/0TZINA181gWZMcF5lHcuT1fy
XfPgeZbHWx2BWqZSI8ZHCIHCaj9tv/kCVtgCCEJiVo2Q9dJ+D+BayOl8TJ+xaTityHvsdILNzY16
zOBgUr1/6zOOfuJlI0Jc5zreu1IrteuXNGHuVYhuh+1hJcb4/vHAvsrLm2rzg0fb5fdsbw0h+HUa
S/0CDBf04MIiwotd+CIWptlY289eSME/Kyq9/JZFl7HGxY64/h+mQ60cNBwNK6QEgPiCia2EXSgI
QEqOzyxmwVNTGpst3KZBzZYEADjTu45GgOekLFTMbVNh0p1hIRnEG60U67d5k3NsJRItCK1hc6iR
TdnWG7QHeQnfHPJhsmjEzgyY3/Wo6m1+1FW3O3rWSrq0t5FdJG99dIV1v0h9s0mEuoQz9W9coD2w
KV/kR70E/7ZRNoIoHsadre1mfklqvVHDgEyPa8dZ5yvZ3+0cXjVPhPe0XQ6E6ToRdCGjfcKTzHOH
/B8mzMLkDrB0uKr3yP4kMJyCwKtE12j/sFZt0nNRWMkb+cAl8rtIfJ1SJsklTgE8bqiD3KwRLOZo
CNQOpRLczjmccq08aQW8qtrrq9ZfBEprqt8GwOGnpJC07SjG/CLxJ5FLJQFG5j05z49k+8BJxDf7
CL7IlfNfgvlX5PZR75E67nueFKqGNSYLW4kK2lcmvWzZQvCOUlPbNLTLLHX2IzieA2At39gVnuT/
J2+iCNM9nuzBifBfRMr1a3o0yaJ+Xf+5iGTk+9PzQglICvPWlr0IY+LTAjT7LbOwVjX4FZ2rUvP4
+5sCkhxRXei/JIEpwAFZBy0/OQz86azDCBDy1BSUAi5FJFGZmWdSVoY7K2kC96KY+hSLccaV/UKw
xcXCS8v9HX4oRwBukjDy37lD6E8j0JAPlO66qprmEkxXOMUVwxO0td0vwpoQp0h76SBNqeYVFaGI
8Qn7tSRJz+77AR5knFO1q1Ut7nrdN3TgwtQA7NI1Muk5vL14VQqUBNYYkLk7SqWgaGogKrSm9YDl
x3rvCMonF5cr+DMq/zERZgcI08Yu+6kiEiAKJhaDZ5ENbVoPKBnYO23vABcwaNRZXCQ3ODc0GID0
927uAbhfue3Zdg+twJE5GS5xJjY8b0mglW+MH7WxUgjYKfUkGSBX1myw2zKqsfXTJp60DYNq+plb
Kr7k4fUeW3P+GxnlaNYFmH4Wk7xJWE0CBaNSrZlNzdf+BA0DnhBoS0ii4EFPoYhWTd9a3BOJIGPf
4nQTmnoYyOCtGdpoRhSWbpDiSk2ENW0DeTahxrdKoxCxIfvh9FYiwNWcnpC2KyvpkBaqBbVnMaKw
YB8WwyJupATr7iWee06c7VTitLDmcEbzjQuaeIsLaPHOdpcrPeNLRqTuiW5BZrG7xJl9ko7mxDqF
RxFH3KX5p0XQSUZguzVDAOAMxVKB9NtQB3D2XvAeCCWaI4DgSp/RZ5mBG3brjHke6NBEM6EZk9fx
qtIuiuS+WPgZTBUzyw9ysPeneHeod8/xvK7iwKbT4MgGbaYbNHBfCiDqAvJ2xfGI88SbYV6AwWXX
e3DrXAi/KMrDem44HWRL5gH4PazeoKTO7QqOnKSz5dJ/oBzWUCHJ96UkWiLhCVWztMrbbqEq3K+S
09zYwIyrzcxIXm5Vf5WRUR9/tClnKuyr+/YGYhp+DiQplKq4Njf3KwgytM+8dD5oYJr4S1xSIBkc
YPuT2Yt2hw6lgkLJOi+irXVZOzzt/JavUChM+qMO7lQmKpM7soqG0b7oKP7CcbCM29QiQE15Wu55
j30/aJsu8/NaSnEXhT62jQS5Zt+e5bc5/JZHyD6+8NjKd+aYa9CjPzAJxhaHlF4NEhb7DXyDxiSK
s7F9iJ9surbZs9kRM8eMlXlSa4Qqo1kHQg1nPN0GIbc4izmIlwoZqxsg7RRg1pY/jKoYjN0P8Ior
XvW3sZGh7askMhMLL+fYFt7rJUoJ6b7bi0INvzK+0Zz8lZPQmvLtDsAnDapmffQSEncwzZRCAjBx
x+BsXOyytnPbmAmHBdFi3e4hlJ5cpcYRGgte7i3SXEHt8Ril9j3KHmAsLhSaOGgKWL9yXiHK4aY7
yZmznSjoeTVFU1Cfy+GI1b5dvs+b4qRpMfZeFl4QgZotPyfHo7lMxwJqxonx/EKJwjgV/0xL3R0j
V8HFIc33AQ/biLCeajHjvwFD7hSZAhcBqJx6JU+d1ltC4H0GaVcpmGcsAvoDUoG77azGoqaEl35u
LNLQIqALz2/NKB62yRHqrlaSFhqHeVrtFWl0wq4GQOv6UXaEwI2XSJhz/WYRbMQagaAgQPBaQX7w
vl6MXd27q7/XrTRHKYezwuvaqmVMyGf4ljOlmP2t0UYIgvAXK+ehjkCE7RXDgfp6bm02j7/FeSm0
mtfStViq19uccLqoPsNDLyZ2wXgrewiUKdlH6VmBDn/Lft9QNFt31IC4M7uD2L9cTz41eJmsLJpk
pvBVJ4A3Rjq5T3IJrAk6c1iJCi0xNE+XhL5tOhZk1Nu6d7NJD5Gvvenw3SQIJUfzdWdnzpC+NbEw
vI/Xo0YEiCktAVasOrWlXXUHhZN1amM2p6/g0LvYbonx1bzXqexBMXwfTb5bGiaVPcANjw2KIOtZ
VE1TGuCaz5U6mvppgMEPvSmKem3L1Z+ipCq/In1PWSdgGoQe7nNEcZfYg0e6IBHUOAnEn92hMicw
hyou56cq/R3lGYjAntHY9hGQQ921i35xS/aeSErBsgaoea17UxDiuLcOokpAfU4evEqgSmi+T6N+
ScHEP1mVIzFMRdD+tr1L0ZGEAibDVCg3nH+mBhdnCKsdWhlbMhOt5sGI1IMA+uj/Qxz79Lfp+VzZ
axqO8/qfMHn/RsXfkt7gWCH/UTbT+5ln686oai2oJ/MKBWvk2fXHCLhgHx/QBDUgpQvd0LtOV7Hd
SHtjPOTtUfwny29K83fNw8ZSGi8Hd4TBBOxmub3xJCyitMzH/gSLn52gbfr+yPpJ5sDUZzWuxxhT
Hf3puAhJ1v7s1Hiw0q2Bikm0kvWnE9rAJ467UTZ/dcyUVyRTmwSUajW3a2tDwETXNi6s9a0ii3te
02/RMhLu917pHFREK4kk4n2LNeH8dE85HW74WGSw8dgECc3/2r+crZmeoo/YkWjASHuwRMHFxC+z
npB5eJiwAP9nw15ibP7AY7ztmr8zqq1RxCNhvYd8jCIxHELKTNxv6rDcs82MzlTtjgaJBRFZasfS
23cnMKMbtqkbRz1qFvCwXwxu69wpqsdxcCnyD6A8nu1LYqX6NiZYTOrV/9eMV7yIY1awGVxlSura
oVsWiGR0VNDYPZVpd8khK64TcPPl/cFKZaHgETZt2hz+KsjLWeWpt3NeObPBeeCwvtLnZgJYxABS
7GvOcYZ0H6FoD5lP0F06vtlQonDqyxaGaIPhXEdF9p7nZyD1pcKs+crWSoj2gWegTTHWko1/alGR
ERhwtdOMPrBsCn3Crw+CKTeHVfDQJwKsITeSIVWooCrRrA6mQud22FCNO/7bDuSOnvJQcV52Z7gt
kDQlRwQ5oh+m4trgt1j6b1RodcBEe4OTweEfc7e59CEkJyooYO3eVDXyCSGZv9VeRiqNEhhfPlcl
5D+hswOfuyPw+j0OOYKRpMKDNC8r2DfYEaASx/QeifR3X+YC47nY9YHxvhHVHPsDxcGmnyEjrq9I
CQbT3LrUicxv4D90HoGV90oPMBrWwl8g6SkSxHpIVpLPWBefKOy1BeyZqkUiYPK3LyyzsHWELUF3
zybwu5MlfPr2LiQ/GmMOe3fIt56r0h+evZm6jvzvbeXvyjck32Sidg3E+2kIiWvG5U/ly/oJEapF
IXbDjBQ7mfRuHh8qh3B8Q61FivMlS3G8Vo215NMmKtBR9lBnTk9pmlkutEDh/phym5l6lyNHOqzp
vuAKT2zO1N/C8SdKbHnibezXLeARBirQN+LVQ1D2I5B9iV7dw6sX1KGaa/bQjyTB39iPGawJlTUE
8SJXhsT+wXCrfe8k15GPdqX+QLm4lToxhriQHKh12IhgcaRg+mhUnqTBTu8G6Nhte+YH1lsgbwD7
P2akSSOeth+2qh/QahmP6wvFAJpAmvGhI8H6vnTLeufIc4n3xcAErWZ0ATEG5MtLJbZG7sTD+L4k
LpyRKJvKoRUJa2S4vIlnZCQj8Rh6T+keXsw69OyXyWj/JisfMMd+yN71Qh4f1SJu0FqSk07249dw
TV7otT57WxcgVfWLvP/6h+VYCA++HlsHGS/T6dEP5zmAvvFWipdS8WK99FOkozHSjw/xUbQgOm3O
SkvhBqFokKevYsbEJS6txay3Yb60OcTZZ2op+/GB4bd6UsqrafK1ARF6usYwjFuw2jhv0/GnP2gR
x4BSJrsMFc/iY83ykri4zl0HqNAv2UsrAaETOJTjAO3ONfJ1ViTf/7iT7EDx7+AxPT68KmAdL26E
xGRZAqEkrP6gDNfPkWMyn+zyc0F9Cp97hYLsMEJMOKfwaR05Dz04bwRaSPW8bQJGFfBzN0RNHRIW
xbceC1GveOn/oSK8IW+krER3KD+ecFpaHhR7xzaZR8KqXkEvGbb4Lgd8D0U8Bnsc82Vty6kTiluA
ICwlTtDITRuvIEYQCxSxFqTActR0ZGusztFXQOTVYCb9IcAF/5pcAoX5aQLwf9jbpKPf7awabsYF
znyOlW4ln6xONRKPOOY0rAZmS+l0Jns0BCNgNfnH6hsbXOQ+L25vzucuZBcHiXWAwy4P5U8SBvrn
9g+SO/JQnvrKPIGBbRWRWNwvhuXLvl3R0y9bn6kcG9eEqyoPeqPS0fyYtn+fnNBs1Wxm6z5Y0O1U
SXaltnQ5XHfne8G29p+6siifO3oUPP3wbE8Kl1otykBo7KF0JoiROeelMewCAEet5FIXY9wBLvyp
kbJi1u97OlpNkqAGt4O4E84DrYxeax7riD/UoEOVcm9YVwk5M5AezFzu74zJGm/iW3KYzoP1F0j4
GaSSq2qQl9NwB4J2bOg21dTeecmbgj1ZEYiupZ/z7n+HH8M75dwhhCldIQlYry5ws5h+RdKI6Lxj
oX1ZSMmAkDnAjflrhmb4Hin43j2cyY73TkHLVOSGnfJ28IWcrxQrjuIuShMNynBQwzn2FjPMvpso
i+YhYfaZpcvsOR89wiujIy8ZUH9WXZl6euxo8yZA1W1gJQ4KTedijWwqzs+HmeDhvd4AFZN7Kwqp
Wf7TZFo+nSl9ju3m8uljVYifUrqw75K5hh1BHGFgwslkZ6/v7FOExuaY35cOo8SxULF5NFTrzHFV
/2WYoYwIbeY44X9DciJGnbbtjcnlPTdfhdUul83ufjcGs1IBOcSa11r+EeZljmtClLLgoedLCV+r
KbjheBFzno7yYPbQgYZzHhALTJKBjvBYX6WWgUszmzTTR3sEYm7gTY0VIDwkwuiH8jgkT/+Os7Yg
uI1YtLvPqF2DBpOV1QPmRFaJ1AtxdmY/f4enoS9AfbrmXYXwv/eNIAVZ6nhr49eMSp3hZv0bTc2R
+EepcrmJ1shf8mUoy4OJBMa3NpSwkiZPEcaUepiZXXqZWyy1GA/+6N1lGH8KGTGyOzWkGWXRvita
s4yYpmNLvLU/4Myj813NTUIGAd6mRrAQYIOTxuHZHZU2wTCHhyBwOAI5ii6XqU61XbOaWyv/4VG7
+7+qIHfTw7LrJuf9+jzc94RkEzt+rT/LOgguftNM2XsP9R+129RCpARvS1k44oMcKa1p7L2KH322
J1EG0OyiRbcliNVABtkZ5FboRZaLVEqUx/fDHYX0l7yig7LexwsmDT88ga/l9aeUodnOK5t9ygEF
aZPbaXlk+OIp5bOUspfakeC1oujNlP2evbx5uZYfg3D5V/h7dE+tbruI1XeqYC2bw7k2Rg+ZLW4v
OIdr2XFSA4vGSXxvDA0umBzAZt7gl/5+wepol4Jwb8VuxVLdDVpF+2WP+3w6Dzvc9xJrnNgQMLSY
L1+qJ4Ezb+rRSAy6wwOUZIF3TaXEdXWqo0s17mrl4DP7axVBQx4X9b3jjuToV682mcOtuwUYOAnE
E8qYLyUlsgU3RsiWENUS3PYPW0iHzwARqmHI6dc+LcpurTMptGcAVTKe5h45zTxa37QQe4siQ/E1
CGv72C7j1Du6s6o8tRFX+LdMlBThQA9uDszRXgTj/V8GxhqsQZgtW1EHKc1aq5+Oq6KGJZkwHjet
to67FJkBo6zZ8DpfGQeCHgUhnYo7hdo4YN6ywH9wDLy/C3qq8pNqQKbPw1KeHqbBbsAyJlRvgpcT
2VcAkmWgdjmlX+/sr1CfcoZGVZvwr5C3f7Aced848C1K/SdNym2E5MjBx071A71u5bFjHXF06zxt
SVudp7wBIu6byL4WWRNt1pQDOxr4OgL4sFFb85gcgHKDXxzMHHN8sl42Cf+6rBfDR4M4xa0eeMO5
/Ta6riNarn9heHILK0AQNilnwle3T167CWgnjsRxEjUe8xgrPzFSxJGpatJSrmrsXHnIb8U2Q51H
vLXbHDNLlzyTwdpOzgYJIlPX4AgAYgDWJEiud7GTrdz2GFInqGzxtEcyjKv8YBly8gxYiz7WiLFV
BbFqm/ktyQn4s13XCMM2cfRhMJN00A6g7wmxMPjUcsVPlMUvGW6TpDW8Z8YOlA+rizCqMV6jSCA0
BbG1YIHAZxx4Yp8zJgxgBY3e8GjgEDzMTydde/CV/pfFXF0DPo5n7IMLNCrWcQPoYqtnc0ItmEAR
EG9avkkFWqdhreHdfnfvcsoLgOADycJMqdcSCfByOhfIHjMSR8AZyL6qfLaOaMWAJUXzMZ708cH8
/psNF4MFsBNPNp5GB7ln2+6zm5iKyEW/KMJAds7riNml8Uecd+TpZ2NWVDiSBiItR/mFoNl8m0Km
0dAu3LTCqnyZpA56mFnv1GXjS1hGjER1nNoZDVllleDalz+b7duelfYv9+tRcKmzvsJPFXHH2BX5
JxwD2WqO5h9b0YTul1VEbAB83lJyNRLFvXdjiPYFUA5UfURFUcc+PVCNYqZDPyjh9dCh8lNqko3Z
SYvqedAzL/aoh8Hwq0hBV+hHgc/asVSAdRI8nKSsDoO/soNahIJavr2cbZlIpr5jtBjzXkcnlbjl
kv7yIRx1E4kdOeE/htVUX4NMOFti8cLBkfGkUHzM8EGNS5nTe0R7hkxniU6nLV/VcMy7A1Z9Mt2R
il4B9PhSN61VV2NoyLgAUQo8xpg//fgpbgKBG/0ABvn1BE4rBSSddIoDFnnXb/ZH1nYK5J86lrI9
n+AUyIayw0C72w+SFCJw0HJ9HV5IN8GkBq5b/Em8Jet2zZlUtSNXIHtYfh05w4TVT7cqZTsrpexp
b+rl1zZdbF3YdrMAzo09e7i0Y6k93vuxreC0eXv/TJE7lMlowDmN7G/fkx70ySO2Ve7ebawfd0RP
JC07Mbaq4Rv2H7w/ivspDyK3o0V/wPAbEvB/jmm59UWUQiETJDAkacolMf2V+CAj1C/27Kdf9ygZ
Vtkecv/CvTOh/k2JMV7MewqzvDooXWex/KthQcQPVR9+MFxQiQJZs8MHflR+10BP7y8z0M5SzIAA
Lfhboh74qvxul/mrx9SKVBy9JNGWr7lTH+Ccam1PsujMZrGVgZnBItsMNs1Ogl6Du033EIu3u5ka
ahClgbNGfBQFg/iQUiCH1ZuyfApcOoKCa9iMFy0eGITzgSNFyVe3frtQEa8c9OsKwke/zYwftdBx
X6AVvarScFRRzgNjGKPiTSTST66rSc/JKRGDbbnR/QFAhUfgxTILURSWqioE5cVtvxL7xZXVteJC
Pe2Z9lhZfAJarrNTxOADXdqao2QE+ysbdX6fo7av4npIJ0KJAeV5lOwtOEPfz/dem4hT6jtyUCOl
GY9e1NCu9hzNtAbA18nWRmWDnnFgGGdKCGss8CKAn90S7bhEhSN2OTnlIuvzDR9HmD/F2tPUKmlM
W/DK1HQLTFNq1fnlqeIIyyF8byOyr0d2SmFbOfbx0iBX5dtfM4FHiPGvC14pIs3yAsVKOZ2NLgYD
rgp8IX0DXLg2BqELAUZLaHQiYLdm7umaU45RD+UY5jZ2Q5YNYOpS+XTpGLjTaCn++XJfrr7xJ0I7
wNtYR8xZWMbrMZAFRJEcX41FtY0abV3v+u9NadpCCNe9XVgjq+Gi357kPpRRv1H7WiVhDDAvNJXo
EC3T6xVQeNnZbJ3XCY5ssoLnXJ8K75bd2YaPZjiGF8jyQLf5NLgeRe58A1t8B43BmkWCuuTxArLo
3F6gwh8Pm4X2RwX5s8HYVjGrRjbStXuiCiZ26/040Jc/2dQZaZrnuwGzHCAgtVecIM5bKvjoaFV7
oAtXi/ZDBXCuisw1B9IWMAo903qiExquKPAqgFwsgsRqYoRnE7Ly8vTAzCD6h5987oml3yuNjDrf
FDKMNuw4SQ06mETr/mFuloZeSk4lYCHXaOKXWfSb3ZU2oZuoqRqo/FF+bxgxZ2gplUatSgSQuDZw
Y09R47Or+04hoMqZFulJpCW73Bp1evG8DOUA96V3w9QnjA9PJ9rhcBcY0GyvkqZTmax8DeNBzn7Q
2GG60kub+dvALX/WWH02TyYVR7Pn5hEHPDi7OG9jCqwVdtL4hOXLPwCtAksJNAFV8xGFC+Y1b33B
EfVOcHUJ/zdmqmcYfD4ViwuXbzGsaoytrf0iNnUkiwxw0Rv4bCRMYVxmjf8Omjih2wLNXtjp2yH5
CoS75xjBrw5Ss3e8vnvLf+wkLFqyS7Z/a7kO+u+pjFL/Fi6r4zt2M3yGSN5IIKV9Aus4gV6E4b9u
dqtM9ONBPxMCKlz3ommNTKKdikGlxYUzSQFeMmUxQ8w/TtwYis/MNMnFstQ2gdNaD7JkZBC7gEUh
gdSChGNyFfawk84sFgxFlW5cY8E37y4HHkdXZY9foY89Bbfc8OSM6V+6r7G8BfNHJGM0+3IBSlhW
f4O5bj5dkM+wzbDRbqTPhgOeEpmhNrTMQ/K3P0BJtR8N+Ei6FGJs2YtFvgADZIQ5IIUOfXBoLCPD
IDzer9VDKV8/rwSxSwfMxS8XqOurDosVn3mYWUFYq8zdDC5hnGm0OKRl4gmDkkXTDzikjT2shvVt
2ReFLBGDR3vfqm0MVlRljM1Vdke2yKR6nhVQkNTLZ9fsQ8Op/z1bofToMmQvM5qL+O4lJa0JCIPH
SUHOEq9eeBYXHKmPBlJ/9XZ16BCNmum0GgAnHvwG9gI6sjrScYzpLsl3VQCaqUJTlZh7cv853sFu
+BICRNUzbO3QxDVe8cQyeD8xrm7dke/+towU3vGV6J7U176vgQbrl1SKps7XFEtGZyruKV3qhC7H
s8HtrhCfL8wS4w+XfirHbOVGqRDAS61ipL5CKcvZ9xeAuceiWcf+ccrVud4KRguMZBKXYl3aWI6h
bK3IdGPTmWw6OvBuXOaF2oU+jKZckesbtY6vYXidNDSSOYHh9iYu1UNP1uSxqrELlFLCxb0q+G74
T8qFLkOxc0mX0PnJz0Lchk2voDNDgYAOUcQnEJpONbvEe4amoPCpemMyn4fMb8ftmzoidsn01V4C
xhwPdgHXbIsoSf/dkaSCtvm12SCu265zerFtOEpdilaNaWqtiCurUvJKHjEt7aV7RS+1zfyT63Zj
M6QDbmQSibF1eT9xTKV/mJWuaKNc3a5cGM5qPiNlZOT4Knebk8DJY+cZqdltwDf4HuRI9rL3SaM/
6H6PhSXJpvmS4MIL5zsZmq4VbB6hovJsKVSKvMiBsRtbBeatoilf5/eqD8ArZ58VUfhuy7S/UjyF
uNtqa5lCRpwhoZQxX+GhKlQjzwtKjcGmR9gNu22i1FLK5JrM3t64rTUOVJrpZxykpnWxL5KLmJsK
km1gQYIk6tQ61Ai74PKLmMprMWNx9RcaE5++0GeApt5XVQaqOxXp1r9xxoNXGB9KjhcXq1E6JmK4
iEzG9eOt7lZNZWN+FggRp8IdQgIRt9sol5gvFdiLGwj8HXSyNmp4FBZp4NdAn+cRIK2pBcLZkdRk
LCpJ8RyFFvaT05EQPPEgB5nIvbx5ofvJFN5jSM+flKIY1g1E0Iq/hsDxigFzK+Xc0wQV1RhJl9nr
3XrRzSXWrTud/j2mK+kiqBXQJMxHL+7R+3I1E/D8euXvncpqQsDgpTSoxq5e0kmsHctO6sNMxa6D
AQ0L0CRPDxCZ8+RjXzYyB2x3k6SiWqRrFQsnLmoXkkZcjxO5S/y5VzWLQQiBAd9I8H9mPF+0tWfw
oqN+B4CSqHWxljsWCMevzPoAKZQ7fKsLj4Dxbvzy6kH3q+mz5VkI98nkwTMYgXpgkktEqnXB0Ppy
tPA+kHoUj7zPIH59t5kzN5YUzJOgs5zT+wwP6LDiQERcSdZ6V7fU7jpxxoTGGXUyYWL93h5Nd/Vc
/AkOcSN4znjZDpecsAAoVWWURN0BwLudgvllQYwEDAGEk2yFtz0r9XqfPOuJl9U+nc+Rjb9ReBVQ
iO/VP/5tBt3R024wR5zNrsgdSbks0Sh7TANFanongG6yvLPDZtMrjqCD8Q/hpBhCbQS3Wt5/L0bR
etpEKxBJg2VfRf/vmxUu4lIoek2ukP3lv1qYF3+DHijGFuzCHv4kFY8USHqEjsFRIgKpx6Gn8HaJ
Z7vpTmkb8kk6I5DZ2/Ya234J7kcztpttZvGCC5PqcyBX3uDZtTa2BzKdQEO26U8PiD4U4Jmc4CNG
nYjhEh+vJ+y4MVgynBKteRWlpe6xdjXJgQXm8ox7aEVzwL+mLjpRcghrXqUJAIEMcKZtmWpjCtsD
mLDV7wLft3NW16NFoAzMC+qLRAdwgQ6i0A9AJ1Tul0vJKGv3ukeMNCwKCpNVTp1mCjh+GCFzCXEX
O38wkSe8+39z5rN1X8pDs0ZrYHMFqNPzSyQXScDqnSzRNLWKsPaT8ggYTjR/p1N2nhkI8gKfbE4W
D038UizbGzYYBLIURaZuuvr2abJi3nXvUXE9TnbAfoiGtNtt88PQSYXVLFh+3gglNZGbOzB0br57
Fc4K2HbI/0ewweeiWvMw8qeML8Y39XfqCfOV3JHUg+OmNsiKg+IBeEckRcNt63080cr+/vWn0/ql
Z3/hFT/K1bt1FhT4ExU4n3nZSKqTUWKRMFiG+0NEUi/jNyYN35FbBai1O08MQRInQsyPUG3t5ggu
FBZWbNtL968F0PURhxeymitlocP1AvdVI1NdqHk4R7ut9rZRrw0umoQ331XH0WP0rWQbgRp8K1II
e17USGLRIFS3ttiajX5ddh+UTL/hj63pJJh4X7mq+sZqtUq+Ngv11T6HRDyS2ZOMNdn85rXxRpXN
vdPSIuTPevwgCGEQmQMifzGPDvvlmHEvu5ngAL14+WygCCAv3sWo3Z1lVn4Ho+55zhnEWVv46Q2t
c0mwgJHhhOcp6cL6PEWsCojTJy3HCAQBCLP/ZbxGqsWadarsbeksjSA0P1HcKrS6JUR8fuhRrE1q
q7yLKu2pf6hV/NgVpbAYOcsdzx8jpHpet2vx4E+i5gGyYz3Kcy7188R1uXiucaUQuKzALbxANps4
MJg0COahz+RwaPjrw/siCxRFkSy/NEIBu/a3ueYdlo8pN/1x7ESFZSeX/mgvFEyFu24JbkSJGbng
aXsyp6UcZb7rgXB+jRI9d6OqeDCeuO5aV6zjfQUatM2xhI2S48RmzUFs9ryv+a3wg0/NfHF3IfMz
wtK7yAigaV9zSKZaynvRHGNlYXFW6q7qr7Ccef5FqdSbHNDTGMMXydf18lOe0cQtJuL9l+G3X72H
GPu4bNWdT76GT2RtHn+LMJmpzY5gyfW7ac9PH/Bh3gXP/pkdM/huJx6cuah3wGEW/F0P3P7OOzlz
bph13RZDAHrNKg4ep5SwtwyD4EVRo8CYWW4yMNXY5O365e8ipkQ5ytFZOyfVuh0Zz+Mlc5sMbduA
D30DD4Blm+9yUdWb8JxWnM00D9kPj6IVG4f68WclO6fHNEesDX7HmjvZ9VE5CnRWryIKKn58v3XU
m3sBLFlp4lpUUgOkSisLRzDzJB3k9e6ou0G3y/01A0gy9sowj/t8/JN9bGm/E7uFUBVz572yNtNO
lWqcjlez3wVv7F3tWecxccn6aeE1xY9UITaeGdsU0Pni0HF3ZdKlG8EwY5i3aTjIzN8NRr7qTvKo
yElOnqohjZDPevPeFneUCXmf7G0T9y1IrO56RKmoXCIXLV14F3ykaY3uAzriXuE3HwNAcRZrxntc
tKRr8hFZtGQi7iTBQP07auG8DnJrWj7+dKDZmXuBRw0viT4gPxKJACiiKdMtBT7cNfrQSvRfH6iA
4wrJ2jq5kaLJ51Ge4ZUBjpCQk0QTVNV+Mwd9GKVM89WfJ4da5iN6/TlMu9p9bwSoPJmjqYiDkZw3
9CyDATCyH1zdsXhLXo5qMG0kiA8AB30F3vpOPe1E8mo36L50CXbNWr9acJDPM7mDePpAzRKidx2R
UqcflkcvcBZ2mA+Dtyn4oIFFYA1eFP83WJyDnmDPPCVhC5Wcx5YeRjdVG85K+NHeCRE3a53wfhJd
wtOAL7sLqKgcT9p9ewjfippbYK4q3ejvfowlJntFJyeVJ6bOofV1zBAFNQtWbRNz4Uh6wbAya4cy
3CSc6FMMS5Xu7uXdTAMlqqy5BXMIEZJ6DDX4xc2AbKme/OM4ruyyc0OE07n84wgkWj6equOfCvUn
2ZhQODv3FzbpTtA3JMxt2TOFUxh2ZoXSVpjp8oIkV6p7V+9DMxCnL9r1VbfS425bV4KXgDVhIXUp
ahkWY9rm28ZsZSZ3WhzTRA0vA4WQVU4kHfaj1yKNc3ULfZyZzkb6J+mewzsJoS8HMO9UDLsIOo1B
DWwIHRjDOSCvpv6IvDXfOT3iXZsyersr/RZj/umQVMUfIg35ihbJTLkpNRbRL1ymg27Mdn9wGiw7
Hdi+SiyQtb05R4wQNznMRgAJhMM0iGWKvNhbpnlAGERWXf+hcx41ccBppQI/mR7SH4m/tugqOnk1
0r2vavyKoyW3Vuqr6d1JF2lutCAygHzWV2v7l4Fa9BJDwJtgsALw6UkBP2jaSGLsfM1ZEitcHi87
D9G4uskTXjrM/EVAkvm9bt04zC85zdCm8EeA5KKXAE3SMvMMZY5hOT7Z1hil9qnXBoHBIwm8Dj3b
yAMkNS7Z1AlfhvuivZBdHZrqlW72CqpYHnWX3SS2Igx2/F2BzvAweLSMY7j9IeDqmn0mhotid9vD
9A7weouLfa4xvCEdtksihYyms6llYxhsOsZwGq2c+X31UqJurqJuk7yw0eFjjNEe7eRefWzQDGxJ
ug95tqgy8qN4RQTVIfaDJoMDwQLRfEKwBz89iBIM0Opoa17G/+XXOST+TRiA+Bw9M5z/eb9e9r3p
KZZ3veCmtT5XwII9w7Afd0zA8ew6yLJ/aRVlBqvS6bBJUxxy7fZHJrLH8hVMI9SpLgvHWhPlZs9Q
DZt0eNHdFtW0n8vRQoNzHhuavBEL4oH0iPF1zBMZQvYQyOoibgIGVwGppwx7gFDxhXpBVRi6I/M9
ya8lAmCTF163taP5ToTdvaa3/fqTtFp+Y9mXFg2TxQml5dreDeNWZpAvSdvAY+gBQ/Ff7Tk9wbzk
zGswuDLdn4qocoXCZtab3N3BZuqKzHo/AXBvE7jwo+T0z8IWFhG9Uzj15CMjJ+GD00322iVGG07G
/dB0R6VYsaYO3Ig0ZQrgBfGNlrA1cENWFUl+iLuMuljlg6HNZnmLkTgr8FgEHsk/wtdIFVaPr6ou
t1VqA4Td+X68d/mtXOWyap2bqljCuGYlYWPCo3yNlrL8yoPVHrPkyBfQ1TytoV6SHy3NoT0DHFUe
7FKgi9TkZgG7RDIqLkUiHKHYETUaMyd39ETxrWEyVyQt94vcbmKXP5G16p2Yr9YExWaOYngVHGPc
1/kOCKB+gTHw1L4go12shnh/xmEKDdSHct6WaTM8Vt7PCrbYa2dzxlfBmXEkuZVUWodWkQ6piZT2
UwzdCJF4R3Cf1eLv3Uxus1bz4GUD/4zrhkHmlEp21MAmXHSf2UPcYlIKHMxVTgDs9NG94vNftpy1
0iseJfao1FAedty3gm9U6yGSjEb8PkiYEDI8M52o0OflmaTN9NRAw9eh0QIMjF3ZT9oxia6Ok/rE
1ct9BwQyKMSKdPZrgaaImeiqeUn/ZAyt1VxNPdP/ljJHMpOrZr2lGdOgnTIgejXfzKEth530YlRu
mwRpOXP517j7IDRInCtWOIgUtebGJnDoBHEKpih/k4a96PW8TjItLGK7KMXCmlNx7whzL4kxwXZA
Gqm5yRo/+7/wiPv9DUCA1YPX9bZEzZjuzVlJRUG010gvdhsERn7CEnlVZIgr4QATV6vrNSndR1zS
j/AF+z+gjPbT+3O/X6P2nkgu6igsN88Q6BEfjPybdjHoHpXP8TlwCDEqpizmUnU+aQj4wLFAlqqk
3AEKOnZhtZJVQn8tt/DHvD+knfDfhGqEUZaluwWGumIDBX/WMGOuuwgt3+YfNHiq1r3BesZc9jqA
hcp96lvSXzpTJYAo8wBOE6wdahhu51BGw7niv1YDuIAkKzHhthhS+kDKxy5H7s7q2Tq5ynk5o80i
Il+Bqza2DAQuKxFrubkSkswjvdYbHUkFPz7OsbPXCgLtC6D9Ji6D9J3lAEdwi8ufPDoRmidFMT/T
OzvOd3oiiH2oT67c+slCb08qw0NMUNn3VKCHE/W/hQj1tIf6xZiSltWrwPwgI1Mm4X/yDlXhxhiA
apyCALhWKl5m3BBC8iEi8tkIFxY9hMivSZ6Gtx0OlPJC8gEZ8gDEFXidi/QN7NTuMrRzc0CyfMKU
HOkZnGR5HKsUH2MfL0GjZh9CWk9z9JUcVsXxGJ5i2bOKuY06fQZLZrmcbKFcsXatHgPEE/x37Vb0
dCH+0z6Ter3yrSPQHdP86HXJQHNlGITwtUCHNseCkU7/dPmYEtZLC5/1gHtjA9DdyDFCnnffdf2w
DnVyDBIYQshMuBaQ3No2fSzsS2cAO9P0hjiMkLdJxeElUSA/UIPwOv/LaP80TqTMItNIMWmS4rqy
5xha9wLZZm6GAJr/jK/cyks2cp5Z7cp95nUx83ksgjoeryrC2bIASIxR+X0u1MZJ2xD1Tdqu/Ytz
jy4LKCn2z99ch5ovtMSvEbm9UbO1V72v/mtfdux9sE5LSjSrethiyBp5iVjsQrlTla+V1EMr/49r
j31wJ9mORlcnezbsqbK+lzIvMYDPJgEounO4cePd7qX/OXq411N+HPjkgT8dnSfxCrkIGGKEGkDi
FX933FsQaKbpeFABEjHXEUDrthCCdTG4KcxepHOmCrhR/ZeDRZidO23aFDfH+gomuvBT0FjyoGCO
gogSfcnmA04j14mXgQzhxP+A6IW353o5OEVqpbwUUrce+4xi39dJP4iW1YAa92dEXLf8XDZ/wZIS
/DMWpT57j3HLMeEPIPuah0DIpgDZGF6itPuO6Ja4SUe+IH+OKTGIq/xHvx7j/+KlfdoR1/AvC+bJ
NFDJIr7JLD7ciI48w0oE9Ru4qlcm7vh4WkniGEk1I0rVk6DYofjy2zNP73vP1PHPDurUkeri+lhx
666wNlC06xBksn2btX6cxBpyXMijGhC8PNin0PKMzohpc3vgiHTf/bVxeny+/qPpIUAD7tdwUWv4
NF2n/eWZUoPbMeBbuAzIOs3GWc743V+xUwHt3PF4MIhWyucs/XXPQdW+4664qJWIkXTWDyztTzXp
/2JbDaxxOx3CVDY3sPVdMFagGspZIrV5JKy+nVWLd6RkC5Ntq8CPGOoqujugj4aAsDAZuRDxiW9a
aHADD8Ddy4XXZL8NcnX2F3AjG/S6dlkzbsKBSFytvnb+/1Sc9zYCx5pTJ9Pz6UeLbCOTZiukcTjh
DLtQfw9r8834RRnm4L0KQ2V/PGgeyo8cNiej6dEnm+SsqzWGKx1DIU2olDob9KHD1Sqre1vm37RL
Tg6ZU5YqqBspb0ygGgK0h2YSkHD/TmBnW8HeMY8kgpPrR59vYUyuKa3+b88TXZqgMD4s7APCgLdB
fQy3PWh8Jep4ZVCCtWPo5LLG8GJS+SAEKHDEunGqIt9vyj4ULr6NLvcNLSlG7+3L4IP0f9TguGZR
KlVU10k/Q/V6uWdx2lUP9LG+q2bDTZE3zs4kty2CR+njor+cUnfBP5lxRtb0UQ/2tmtNB4hbsBJl
cZateNkJzcwZ3JazhB7Hlg6wJ8IX37J2LVz9+mCFfTaMBQArQG4mXm8hyjyLUV+9pJhjhUiHpedV
dox6E9XnLaAj9e3v4qVRgp1WVrZv2zYkSMmo76Pt1v1GVTIRyUvCEeNXqvmTMUPKU2/e5WV4cWxh
ZzF4tRN6Mg8gDeorhn6F+irRxQ+kyYB3PNEMqSBiYS7/5SzhG6Wu062WgTtL61ZCh+85f0I7JUhU
AXEnslUNKxXMhmR33LtCP+L98oiGNBlolp3lxBbZnMBiKujqquFdSXMnFLckNRhltRu4MlfE6UCv
SGw6o4S+4fpGsfZJgy6UnGWNauSJma2DF01izjE26VgZ7KaIrhqwbei3zWaL3JqZZkH0P7LjPqvq
FkgHhP4N8qp0Kvl0hMM9nwmAC1salh/75zRXIPZ6IzAxY7X+MwwaVgN1Z3bW5Qnf2a/3W2YH2MwO
8pF9QaKkexhGTO1AoTGW/a5p5Ige+poRiYwWMo93wJ2F04n4NCrtXXDZ0aFPqjwwMT6i78sl4AKO
2H8FgxzhqoGxDwmG/yx0ZKofb4lYpGrgIslkydLyHc58OoMsKSgIurge4q/P540/74Wf8OgFkdII
DsjeKd7weR4GfjtCY7JDYlDJ2KMcrUY/vsnguCUidZn5dvX3opXWCV5fnACQE/bjVD1NnQsZ9YoQ
V6zwB9Ht0GGw+uHGp1fuUZ29iDhAv12xFyWuX3qfHN+4+zoiyOK2RXQ9kSgw1dcMlRtbUt5Ryt+j
C1D6m5EJPKJrhX+L7+dKvwQdUyNQIjMTgB9zlPf1ZyMRdBEC1qidewn2Mrcdi+1UbYcS+XaTBCRb
6GRRr9bGqdWrSZR/HrCeUY1tqJ+V0P2zAI6PVlwBNn0k1jQx//pI6rm88aqFnVkLeDWO0yLL0xXU
Jnm+6BI9W0R5wvjoh3Wx9iV6ErFTsCGeojSa51oZSm/sTspZkNu/e/ED4WhElD5zApd0AmA8Y7m5
pPiRu5QNJoF/qCRkRZH/i3bHN0BGhuJum0Eunb8/lWQaW9XJOE3izhLzWgiEkQFDTKvtXJ6tCK9v
A+cP5ngel6ncXrn0rQiCfdQaI3AZCUCOv6uVI7kVMtTtHXfBObVcySemohTRM5z6/HruXqVsfSxO
5kCl+/eBzohafjwa3bjdvKj1HXt/Lu+yK6ftxvr5ZfUm6R3pHIy4TztqQnkRZxjfAIbWIeCcUFkN
hnwYv+541JLlLWSE4sMJAmzNBYqh7moqEelfg/RWqrnyHZ+nyUPPiF/KKiOl7lSOzFC4yhD0WhG5
+XW3ESF6pFIcNXryyK62LH0c5mnp4ophXlWN9t0AxW79o3gaCbTOZHMgPCh6GGl4pW6+C9TLuD/F
kZUlolvo1Bst9DqhBmXUskxXEUmKgpuKTHSwUM1VZ8YdR6UAzIEJMMazU6wJ5SYYp8Nt8bABAG4C
/V3NnxikSLyLQB5W3U0pe3VlZRQZM0YIOQJO3SKpN8xuWbq/nAHLAIrZ9uE9nW7k1KxfBneWIJo6
KZBcfdw7HvENH8Bls86xX+al6vV5yKNz+LcsVvudmldi0BIg2UzleZj4vRmuU5tKVEF75dXu7MDI
68fBbae9DVtwg1GD3Tn7Fde4LsC0FbPhe1KUwZaPYrqyxPbsGK42AWKJQbVnHxCXRl+RAk563kz9
8xYHj45eKECrDTJRTqiXcYQUAaY4SPwGkIm+9TcvVG63tdefuTR3LNcvE2N+NMez69WcGrkjIVo+
0LtdT4Kshx4Bk9HSHJ2BDZQodX7U30FtxvYjCmbP7R0zZEsi8kMaeFVtVFf/p5unF4Wv+nqWHKdp
Sr7kp99v/4i7mRiqkXZ+0N2HqxJGjXyf1DkhrqjLedN99GHHlICL7rZSQM/sj1pf/+bCK+JVKRsj
KV0jrKdN8Z1rk/xLJpiWZNtg+GFgkxLo4UG4ETe2WMQ02vQIb39yBd6x2iIg75RmAzDzRdfAfq3Z
aFJzDKoh20q706ia0m7SZ9LBfGXO/FCkQTxeCB0hCNCRhOjRSUklf9OAdQbOtBafaYlTiZPedhTg
HcNX0EDpq4w0EV5Hj4baoSHd+xnzmk7oSohKtw4Cbuw/sWumXXpkWjWSxMzj/X5dUjjkwe8aRpjK
rjM8DzbLuJmyaAQcYltq4RmK9CEZY6ZjaHszfnAfOOyRd77USElG0tLplMDKEgIvQzcoJZ1t42DO
J8pLLMqEcfaojKK6/f0+4QPgJOkUKx86PZOgd3Zs0DA8EEXvvYsEmx9IGMeIGXtewiy0ps1JhPvS
tr5SpOyxtt0ty/TpCnu1+uCpzxBYqPR14iEOZE+9ajhq5cgOkTKGV+TUSrBY/GkSOE2hZHaDspDD
K6dC/toQP8En+zYyAuPij9dm7boCIZ+uqKUts7pe50/vNOKaNKz2renclpMNDy+mZlzDNTYoVhsF
uc3t5MjUGDlP0bQHcWz+Pnp73IL6MupPDukUxpNKwBY9GTf/QlG1MM+HRft0P6QEiUSrIqllFD0G
4fz0riNA8vSGaE0ASRLIz958lv3kAyRIlRtKihnu4kGyF7nZruBVGMxBiKgwO7wwJ5d7//pZ/NJ0
5siR6Bvy/U0brjL4s48HhbNadzRf4XP0tNxFe8y1uc6J7o2A4Rz+Iqivd7REMAqgJ978XMupQsM6
28eDQ7dvM6o7cUZTR1nocGgXv4A6O1vrCDPjj6xuhMoSNSqkIlzewEMTL5bPNXijaqYjibUT8tNg
moZR8Cwu8rOk8n3k7kd5hxfP44/IuopgI3War8Gu9FNLceVZgVp0FMk9kyZj7wogj5nmAHfxllcl
DJ+Zrde4Um9cYGxWpFJuXaN9474NKkkRCY+HRmcaYSLuwSSWuJT4BzYNcgDKspS7dmodaShaCtvB
QzFCgJUxtU7fHpwUHCWT19iE4RnHxo/E5Si63Q2eDa5WWD17O1/9NjFfyktxL81qTyLkeZGkHorM
KaJewJX4HRn6l+1ORLUjdQZfontVR4aOJgxyGwOiUKnbg00hNv4JYpdQcK2NaBrq6rDVqRQ4+lSK
sKTzw154Ds9xzrOFGUwkSjc2PY7nslyBxx+Fo0IUrTkhJiEkngWNQ/TF2n2y5sR1GNsu5nYLroBJ
Cq++AUoE9bZq0E9TSNtAEW5DRSUNf4FE9ZJRMICK5PqZFwp+KqfnCCxZgaQJ7OQEJKhGZXVh3Txb
t4PzpDQ0yav4R4WMDKMndgdDi8OdgRYaz65TC5wuiQFnGz1UsHJcw4uf2F8jrrdOlln4U1/OB3qW
U7mDBJK+4/iFUPw204awDktRzqQn/wUGwGpzFIczgjYgny3h7G7V4yXtqM2nx4ADlTg2lcAvCRDi
H8I2tWq8CwheYJczV71QjxxDj+veE+84c2BO/PmnBitWLw+2uBOFSAZTbHt5mCBDs8A+j0IYFMPG
Q1ENnVQAC9ebSW+9RjZXSbWi9nQm1ZplCsnvwL+0T4G4mGdofosZj7gwC34HB1F1qRCJzyJFOc6g
wuxB1pmFX6UR2bdJrVR+uCfx/swl0EX6ecmJZOdJo+ZRdlXmKv3F5FjFCTRpRK8kTsRN2j3FEiAS
zlZz/m8IkOdwdCsqWclnfz6u7sLskYqMcXfUtBRtGjO4wT3Lau+bSLlPjuX26FcmAJ/Bkfq1flkB
WnNkJjWCsbLjMSPZMp0yIFrmYyFdQWUQl5JQs7ggjBSVTAuBkaCTzEKAJkBM3Oyb1lWfdwlAexbG
UyH+l+Z2hFVaVV7BF6VV0zgZLvjMlEl/YuHrnNiDYHW8AKdT7f7Saybuby2+Xj4a8c7kq0zIQ2lo
qpq1k2DJyx4zb1tMn3IPVbnhxFrYQGgrdG5X7EgtHs9uEzSjBTRDbLe4Q0B31JcoLUAcX4mmXeFm
9r2PSc7xMKgR0cVleI/LgnpCuYUDV/kMZZTf0iXOtS5DnNKJyR/K5elL+14p68MMtuLNA7Sn98fs
5vzM5O/lKIC6eWg/mssUKMAxrEQgqVvLjxLn8agV3htRlRJUz4Ntm/WobDHJThh7GQ73LlVRkYfu
T+Xjh7aD1jYzE1hxOsyokzfpJFYyDC5KPWOy0jN4yanMflaluIG/zpfvOYss2ZBmpbPsl/x4uMPP
+lFU7b1I2OoGmYuuBWi64eqNzXqXZhEC/4As3TLZM9Yzia8Fs4Pc0h5Aaf+nesHJgxQtyOVvBROa
s8QbRNLXTdZeb6OOHu7shIWQ37G9YBOMgN/pQikrh/kLCfhgla9+rhrbp1qAarbgqR2IlNxZSyD4
kHqXT02TQc1rpxOdLqtYPtu5s3hj8jGWxe3d0E8wA6DRkieQZ1mzx5cN9OOuQ+TwiwHg3PEcG1JM
t06z2MiTgsMGZWDPadTdG912Bz+FRSd/Z/tr3BmB+gIhT63zQwm+lIhrkEld+gyQWjrVlYxKDi5c
OkKVN0cnuSb8w5cbq2X8Q7hWSF+aqIL160O3gMrBWVzu5t+og5+uktzv8MRS7CRCt/DPwuk0qSs0
xNoBlI8LD2q4xvKTSBOWPQa2LsZ7/6TxcOWcFe5g+ZMe/Wig0+4BoaoFvIeC9L4fWwtgjfVFBkLo
Ez5BkBcLRyCfbm4CCc44+zoqlKofbN+oYTI9OpEY0eoSCfjziqnsTzGYpYSIC2f87vJqsa7iNwxN
oVMrpEmUf194TsZHgkMWvgroJctCOj/fDzqcrHZDeuhTB8L+G8/GPpQeht52OxzYLS6E3E4vSmcM
rv1njSlyEFE1v7PwdVN2VTIhryfM5EVTS42YKF1WWcq32yYY0xnKU5cjFp3rn2S1xmzEgcs+iK9F
i3j/W4xgVCZ/lL0n9n1mIwRZCuPTAahnvFnSgW7xOxM68+EVFN84EYhVW1Ch3rdaxKS0ZhKdFk+s
LRupV0KPnv9kpVKPjE95xLnL9R5W26oTqBjsu5tkgQ/aT/7MBdI3PfPyrORAmsrYSimbyMgemdhc
TbutSX5hKt6ExfaQcSAnDMMPPHDwY4jsuNQPP8pHtQXWBbst+F9eqXX2wrveBppedQzDH8GZc6/V
x30tXtM91sNXuEDlcSY6Lsp2IoWsveKSLVvOjen7Nfpuprx9yT8GOXu6hiWyYE4+pLbZNqghNuRy
fFU197c0uwxDWuVE11taUdoHbW3MhwItSoWZZSG1Cfr8PdwU4U6WdkrY71tmtrr6l4bdbyuC9vzl
3S5vM+VgMqA5FBkngrMX8q1d3Rq/dAfih74YiETsQ8cYO8E2TZBXMWOTvs+SFyWIc3/pRoendrxi
BrKJhODnuE4Qt+/96VVxx73PzdVF5H3RaFpmlt/wBW/FCLNJu5oSNwX65BgJ4XybJ27oNoOWmv62
8i8GR9DvkB08XUG327/9lbIRc9MPeTgnsAsPFjxtHiA4NAoZmeS/r6Pkim1eYEkUebcYA2AJDoDD
65XR9oatAB9x3tHw3AqQTAJaNKZ8i/PCorZaXF+qujB/d+2ykyRJIFg4bFK6F05Dao4aMCoy8zsx
XSx9b4G5iIeQJ6mzOHEVwPrilgfu3rouSePKJVGEVEz3WSxlljxttpA2BcF4tVX8sTQeiRsyzTvI
m8/CdDZsRg1/g8j2fGhD6d9Ut6KqGwI22RqlAIE6PTDTwZjuWxvuHdp4x0YfuHC7GUl22mlyBi8G
Kf1yRHssgc6aCAJzHQzNhlFlOhrjyWOGYmmIIK29QvrB8+CHNus7qM20m5ydPEEQQNkYL7EC2/xO
NX2YnD2HHy35jHcn3ysQMRo9IpSvdVdOSFglUnPaXTrsGTapJ2bn/oEqFEIfwydPS+2WTuy0F0hZ
aPv4m28rBmPEuDNcz1Aazt5Zu6l7YoBHVYf2zGUkYQRYMQCqbYNbHVNwkxQSfq4KLEAeiYeY7Nwt
zWi4PkxDtu9GmVQ8er2JFfMHeko7XVBjFs/i4qR2euvkuahCjZGF40xf5ljkQXHmRHBnyupDHsgw
VzMe7xS8/SRZuuM/98fUMHt2jq7HJ1GqLtPTcqIXljH/54CX4Zw0xs7gdrZFi0jDKZMkMH51p5wi
eohRbUhOXgAC2y4oXk9piAYjOqF4Z2Wxtqzb1Y0V/f0dTLfyBosxNbGrAbDbmY7U2N71zwtA7e6g
noXxs8T7TFIvGediVJvphR5cgkV86jtThUwfRNXabHIDcBZI1QEYA3tYo+B+iXIZ8d7jdEOpD116
EoR0JRSB696dwpxIoo8DKroEKkWHiFh6TFR64LSkJSLBjzw+7UWNpMCvE2niwXqfWrbiqeqhwSJv
8YpMFlsvRbDhgOOojUFU9PBWaFX8tOjyHZABmn5T3Gt01TCP59QZkQYshUa6C6VIe2Wum7Md+mSD
q2Jz9hz0P883oUa6Dt+Bx+J4xeyQKirrUGMslc1+0NWRbR0slE4BnXTy7mkYi+Li+QYHJ1/ZW0D8
Lat2f/bPJcWZ/iQTlZhmfF0BwxBIDQKT0odzHJ3g68Yc92Dt0CD2wR2MyLYnUclZ7gK4aetUzVHd
3PLgxggZkw/kdqpBaAf7FlS2+YZhiJ+rL1tM6I2r4V6VfwZmtxdFY0Hx1cLuNprnr/6Ol0OXzrrM
usfvS4UnpnCEasa5o+mNqUm7j+ehAC0HLkHfWwjXpou+icqF2EJvrK2CbXRQuzQcBPo/0zMurXbG
Ocn52xOFEIat4OhoOo8XhlRA6ekZML5KtwXKEW1mN2zMtRs+ZL6EqEJ1WKS5PEDnyq9OvRnvk7bz
TncjxPZ13STqtlKB4kKICjwrtzwMeSykYXMIKy0nnSPVoqF8ZEYov6+nYRwvXd/qW4229XlybWqk
11DdGtDJgHPsWwneqISBF/Z1zoo8oz7+Kbj+UUCjlLZcaq2rwquF/CIxHzxQw1teEWdbUNsEj/Dr
ugKczW1QTOVPef3/d+jf3PupdufwCBNZwYbWEpyeW9yzxvQeW5RqAEjw99VEOCC8n7Oif0rB0wHT
CCVKBJimiR7YrL+4CmtjOUrLqvHJ1jw6n0QrPUi2DKX64FcXMLA21elRqEjkr/5qEzp/71HxceMh
3B9B8MRUwm0HZTbRHGFVuqgCSNV/tRpj/vG3GYNzAgV8Vu42hzyzRavL1y5arOhwxAFvtVHo1MhR
S3wbKtpVp9tSXODGX8K/2Cutlv3ykZCKbQVx/nF41pP8EsR8VhIQiRdPn5lH0NTuxo4hOj9ChbIs
nIwD5y4n5sEVreb9Jz822tdOcYvpRGx/kh6r4+W/9gakhA6tApbzZuM7lmYUfeCJBCk24jB1BvsU
zddquLvjGs29VE34wLBofANCA19MgOLlCXHx609ZymLKM24I33Zm7zQLOBmZnoktdYwG8Cj8CGNj
20fN9PHIfNmxARPA6Rbq7hJ82qKYzKrSXjlRfT53V2ffLiJcU/yzJIB15cIUrJSi2Z6M1qfXT7dB
yZvnUi8NpMnpeU3d7lDDFU4pE2rvUAKUGK7yN8RYWWlhltFXO5bIGLTUgnOjxS6/LbPN+5wczhOO
RBEqOY7UApvBkeo9ZSCF1ZeMPv+fSgxRzS0vMu/lHw8sckkfKml6DcLz5Qzdah3gcyss1JcdCORq
sBEoiIW/CaGbINfFvvbxYK6JXVKUvltsujbeSjdCKH4yHlucJ8j3Wkxt25FvcSJXw5HnGf3/z703
nHc3+C0jAM8NT2T4jRMveCB4+E7EPDnijBtzU8iW3Bzn9I9sj1hVUl4KDDkWS6zNxvAz6apIstpj
AiXRsdU7PB77HbmtY0obdUhU1tELXYz02WtXrtR0BlUAhqQFUNtCb6xTMF6ignrvYB92jJF+3nfM
8qt4eNb4hLy8SX1gxejkOxYeyZtRCsqMzAqb/RJhEIEBmWMg4NKIXONCOwhrnImKmrRpb3Z1NF0u
IiGj3ALMdgwFKGO4g7GRmy+kZXHXjzU6SzguwWFiaC8awUG5vL20qHNfVXPw8LdS7VVpVZ1YTG5u
x8dnNMOd3WZ06mRh2ILedEKAwyWvLxWFKr7giX2BvLRCWqn2yziyt4HWMfJALoGdacEr2HJYSBSv
R8JpYL7D7HxWKpGOoWrdp4cxxb1aZL60CR/nUlcGTpuOwl5LK3lFregKleZTHYtf/EEXxmkpjd8t
4QuMhyQeT9B/aXzJZhCvrBcYWlz1+jZ5oASBWsUKFQHF8Fj8dZ8AGLcLbZG9/krZxTqD5tuD6he9
y2WqCZjR9GfDaijuqXC+9hEzKLS5ri/gw4wkMjBHSXv7XgTulGgiFkkJtzOMWzcAeQo2Z0GBrWyF
PC8AEqAchIoip3azmwUtJ0JzoB//zPbk+wmJvvPWpytboVYJmov4sxSYbo5zmu4FsHVEBC2qqI5Y
6QoRiHt6hS/JvQu7yX6UUrAr+BGKI2tJD3S54wRONMjtb7KyeWSYmla7Pyh8xOckqE6zrxAjkTH/
1MOuKqPgHUAg5fGNu16zR5Oll1a2FUzA56eqFAyW7tU4elktM291weAtI04Xb5CAwFZNXEka3eJZ
3jhmR3XReMI3EERl2D98fY7ALzYk3zmiAhGG1DEtpo2mB0wrF4qRS+LmZypCyZSqVZHYRAcNO1HZ
1226b99mbDunzCa7p9LEtLfL11wNA2yq/dSuCKH6PvOhQVm09iUjD+KqR1/iDSxx+pl8yhAOevAc
iOSDrluOHQZVICKwN6dx/zM1lWIWQPmzB4Oj+r4HaOHDqL8Trr5IfLlWFGYVHWVM2qORRW7/Krxl
JWDXazkKgNI3PsKss1amxuUTzWCl+Bx6yUOsNBHZJU0xQgb0LJdD+nOohVVczbDbgQY3yTisxd3/
EYtRKzxIoo7anncakKxDxTMjEBt1Me6qTticG+LeVVB+/jeSLEJcPY3QIqAuu0xTGzekGg2DDPC1
09+KKLQbxPBhNpOg7GnUNQG2OZOTJNppQxldQ0bm75jOwKMbzU1u9+CNQKTX2sY5SQ0Q6duN8G//
58VHQKMWjeSSj66ceFFFbsLu/bCzAFUe8jcfdBtUsYB8k6lwwCPLTZeAdH1PPH99iunvoDwH+GmM
fvb5XegVBlkRMpMMgKj6xV9KV3RPH9R2hxBoUXYJq5EiPzdJBp6AVkwphQsxooea4Fd0gH/PNR+d
6XRPjK4z4iTLN0JK9qXmMJqMOy044cp/lDE5zmQChnMq5W13Wa+Iq7hJe2T9NN1luaJE/iE14XZ9
FQumbpCI0JAElU4bqV3O/hz2IihyzPH2E7pufGEB8IfRy+tMU3OtE3xL/TFDovKrkpaJbGqN1c9d
DhYYkjwsiudZVoZJRvDshNh7yZudK8AhZgD6CTLLKPSpq0cW4J4ARtASzPx1G1kRdjymS9yl0KvE
81//tGrTQulaG93xT9saPRILvY4W35p6ZKm0JLK0Pi/6UQFIy7Ae5T9MQzIgjQnxceMgN145xZgX
iTMbCmO9OmIpcXmCVldtuEWsTPMwvwpjkgJ8ar1fnX6tANAd+dZMI/bZC0uouoINnGof8YYsUiBj
9DJ8yMAPhWCUVTTKlwu3gFuv3ARREFl1SJXkvWZFAYjVuC6xI1Fn2MAlz3+VQIpknbLABLWfOP+V
g3NXOe8wXZNlbHSH5AtLLW+jqPAhMN9tywW6GINy5IN3DWwi+lsZ+gHoDIxYd6FmAFXhg4TieLnP
oxsNKgp11cBsO5dnUfrmR4lIjPfxh74T9OmOKK7/3IOHdlsrH5EZLXanMa34vBEAHW/5+4t8CWmY
+O5avWC8+nPpP/eQWKnfaO2LWPosHs2WH9Sn0CC1F8pJdi3rLJcjv2ETTJFe3kJuHJeAaeH9SgFu
ZB/NgxvCywN4p4Y5yjekGpNwFCmdDPoVdXh14QtymX8Sfev1BLtPiJuNxr+ZFLbSfflpoo9FAQ/e
YsQMvKYWXvCjf1lZm5pHZJ+gmP6PUthPcnIOvPEhhPyPMNdMA4fAvoWb2QMjEisUsFrYO0oNbyEn
tI3mqesa9sxGNU8pJbbBH8dI14u6tKYmXC/9AqjNCLk/VO0jJ2HXyJg1EPQAOjrP/94oXTFoDsBA
L6m8udrRg4DQIjbwvgOmKXsaNFHWjb7P/PDgxRM/FRCw2uF0hWdrDj7De0oVQl/ZfmaBZepX7OAT
mKdhR8Jzt0RB3jPUotmYJVs/ktPv5qjNQd/JsgzxEI0+pYclZjXDtP8YFcfBlL5Dms9xn0NoRJCY
/nz7K/kudf2Wxf+zE+1fm3+mdRI9FYJnZAcoAcPv//xtTLTDnXPRLvDKaj0f1mCi7xaRiMMV3kTq
NthMSHV/+HTrKLZ+35dSL/0i2W895amw2SSPWz5QzhxgghSQsPOsQgOjYH/c3vIWEUQT5tz7NTgD
DVoFCDcBBjDXE9wX29rZUHmxfgqFlxPc4E2EhI1UJfsUQTGHfNhv3QXBE0c7wM5hxOTY4uHOTqhN
f3ffxizsFPhjoeUWNTZqdqXyYx6KE8cYDzdDExhyiURI1ipJhhLbiEhHC4nnfEag9/pKSuEoTdIR
u8TfdYksLswhBZ3qzh9oklneArwiZ6QzIUk0Rb4mKccmGfNbKbKcGlO8c6WOJRDDZFVt5+eEdnwQ
ua9XyIpYzyM64yfuYYm+CLQrMdzlWs4qeCX16NLfPxITY7niZnvsNbiW4Yu0y7dzmbvxFo8juFRR
UT+LZR1QV/yWWldR/rKrj61F43M7VUxx+6ETAwXIz03/0e7F9TJZEjvyvCfyGowuw3a1NedKbQBE
/LmmMTLatGIRs42EZUCF1iidDBLNcE4JY1NiUW2mq/kDRdMPT/ZwW+BE0eKanqq1AFFpzcK7uRGF
SFpuxF66V3ntYTU0APgfY6OBQDBRhIjwXEgXOgVzT+u21/mPoBXreLMsndB6kF1KYQAgDVuN2afp
XT+0oB8fFIhs0/JoRlkVctvyIcvgZiHmbIt3cz+Gtm+5CSz8SNA/rzpHX5ImACDnmdK1imJYgHm+
GMOU7eV/R4d7C/1IwkbUAI+ftdvaYuJ4RsoVCvlm4nEhr1ztH1Tne0eA/bF3kBSbpFmXypa/xfVX
4JQodU17w0vbTEIQXH0eVzKSO7kDJDdQloXySsStDvcq4Uhw8sI/re/2iuv9+VJiTDe5/csBlsql
hDAG/PdUnug9VQCgZz0LLK1fKos4nXn1Xli1u3MVe0tFW0xNSheAVljwK6T1+FI2xb3MNX8QU4rP
Fkyvyasbi7vnkYhYtjRHntk4maxdJzyE80y2fPg2WwbgrxanXk1fKmcZUKZChbQz7EBeI8wzihpL
1N+8hqoZ9WPGYZEarApCszySxY5lhBrXgJdhksMdppXvrmYLpRdLiX8P/ayTiFZ6dMySvFPP2xFj
igMQvESIQLsMWPbn6Qiw68FRPHQh8GadGgXyKKYzYgSIFx/JGGABwyujLxl9h8tmb3dSisKkdLi8
azlJwc9tZUz1u/mFIJ/vORCistCBLg5rFvxGlMrtJVBFGmHC6dT6M8EzksesXtdTxY9sMo+4z+m3
414y9HoNW6+M8XcCLYp6J//Glxw0aIIjq3OXEgjcQz5nifFovBxiWrWvYK9ChS5WfSG1v3NIKmsF
sWFiZ/qiGTaH4JkghkmNGeKvM3S2/SPFCacej3GtmCWhd+G+DaOROt+DrbYPFqbmq8jBg5pEL+0d
+7/hYu2T6IchEFWsSVRBAtApmCT/72mnFHEu+4aUSi36WWMCJhYpu5X4pnjbNf0q96LmzWaWHtJ6
VR48nZcdAn8Yf0nnWJiROS531h7SjVqXFjoeGdCnV/nys+mhORNlQlNJr2izKaz8ixH9mTpFhiWF
HF0utGzm8tkWd/mOph0NUD9YlClhGLlK8Q4XxdU5PgQyuKTUhCS75rGvn9RMR2fn0AaDAWrb/swZ
ExQBQ6WvHd3R6iZkCcexJX4F2ByXBZu6ZfzXNkjateRHyqQajr/B7Ts54OfLL66E6LFX/Evej35n
7t1wzZCBF3X/2xGW8AacCwd4eUJDgTlhN5NqMvD39IsBvZbPu0DC7t8nu9sck3BEKrB2fpzZAF4r
7nU2ASTbhbvj4jqiP37tJwHK9JUjfFDAM0QvwvB+r67oA2+J3ELGadtrqMUSdsUJB6yXHcuCMSWC
1IZQNECaXjMzrU0AKrO9SxNAUnzJt1ij1nHVwa6RAtBTHP7jx+MzvgRaqFlAJl96wU8XD5xnAUep
CzsCoBF1sMSdI/GWLTPmQKYya1JJp7SyXTAxNXZIxpw4IMAvG+5694pTOvKizxazrEscTOEmnUhi
cd/hGFai/SBa4cTP6IJ8bTaNVvVrp3ynGG/iHAa3hmMYJddN0R8sYudHhg9c9JJexgsLMKNM3UHY
q3SpRP5CpoNVzGz1YNkzDsGk7M3On2l21P/iN/usi9/DlFAy0CiWlkLKGcHGbbxjG9+ci7yKMQSW
MQGnz2BE09jO+sopCKHxmWsvJuhffoA2/ZQ/IXekzMG+3ekkVaobEJ2X2Wf3IUm1uy+0jWle8/Kb
Ukzi5JYvaZdgSt83xq77ZayJmoH3qbf942/lFTMhReHbjvRGZQ6RG+SDI43+fnoh4mUF0UiBjtro
W2OhG0PnDNAKRpspjB9BGAFw7VrdzSzyPJxwdpSAD581eNqi0PlRK2i4zcoFVTIgULd1X63VpMFg
HNuEO21CxQDDFZpj0bK2/1Zucuda8+JR5S9KxlmRfZjpe8SQmdZWwBkKQdLJxDM6a43pVanwZ3zJ
lqg8ROVYN8VtBvuUQ0rXp/zYXycn40E2w/fZJ08t82AHrWEU+zIDnaRAga+v4DqwJf4ZMzVnnjZV
4edBTjh4wzQUArG+waP86WGZe79LM22Wd4LeutiR8aowtqBPZFy8mUrIO47MxOYlD4u2RA1uoL2q
dyEh2i1saE1Eciiy3v0mWlXEH6c5w54p20P6SBksBKviVv/EJzVH3hb7od9BRSaVvlGEYLTwE6oa
TxOXqK8sNWqO/JVT+Q7Xh7J8J0V6inFR8jkY50+6XhlLPWiZSAmaS7spMGlB0Wb6NQ6RG/3L/hS+
5hCDvllt+1bQ/CDi8QVt9Uo4tebBLjzNyF+YyLMgN6s7WXedtA3n/XSm/9lV1ABs8dNAY/gadj1X
vxTwmclyNLAmBKVVQevg7MVCVhsHCAyJw1xSZcP+zBW0UNNoZNTJ/KRZtTsTusFZMViabRqJglDT
HT1jdmSHwKL3Ow+QMY4yTI6KA5lUUSWMo33q5auBoiWNuawnorNZn4BXaqGd7BUS2dSPZNxnVnff
9hcawJDe5lqwtUkCsXymW9Z4qCYv8wpkHOv3CxGbj22ud9/jqsiNh0z+bgLmftP6Fv1ktxWWoEJn
9Y6V1NeypHCNu0t2xixm+zU62RcHfHZA50Z98gj7Tb6lvUcslrZixF+wuw1Gr0ULBcukWqsbcIfw
AHN63SAHM3KvrhcqwwMXbacApOwhkTDccFOPPNVpzcqKfHGKHlWjhacGpu2G28bYJDK2CW5Yhn0P
Uk5AxJGKH7OYekM+2Exby+yecL+Dt6n9hqkFZD5md++SthlTWB8CHXRIFfI3Pn4+axAhLCnZh0iN
VU8x7tnZ10hxuiKwKiuPVvaGZZLvN0LPK+Q8dsbIQQ5WRQUjhl1IIf+yYWCOBUvfWW5OSEwiRFz8
RbL44Ua4qOAdn92T/S35ZtxMp2eHQwIlaeNoGLNH39F6XBZNhlB/bx0411oe3hDvQe0I8wO17c+R
e+AdIhxgkryJtXHF1G4cAyBXOkj4PzFKnNRCymDKabFu8K284qIgEPTUmJ38ZW/2Rkcgookcf5l+
bigq9gXduIAmt5lqhlFmrYb1XQcEM6zLLdKNQZWbNNkgsYxsWOl/3CzzHajsSMDCLLjPqWFoD7Ly
HNT+BTIRFV4dWHAeTKn54oWlDGaIZ2KRvRfNzyBfD6wGBhNjhbDDxSvsZA/lyC+uF2BnAYVIEpRd
3igWGs71rnIIvPoPdW9E/LV/CGQYIivv8Jl8L0WkfnKb5aNi5dUCqp61nscHz9Gamx1ZOoZojUP6
nEUCMBEqu14heWD7QZl/yZqAUZPSsJ1WvuXDnlVp9vTWrMOp+p0WendueaqEZdM5YXxisUmpPUup
8iaQCE2XVuqR2t0mDHSAidFw7GDz38pboj8hn4JqlRoMfvuCAW5zex48T/JPyZ7kpoUVcK54lwC4
I2uKT/s4EH85zHdTygIN0TywzIt1EwKf+w7fB1gWKNEbf0+jW0gHXI7vkR51LGVC3v8NuW9W01y5
In4liT9ZECN+brUwSh4Us1wuipJr+VCbykKaXhWqjySYs2lTZBRnhgj/UVGvHhObk43ZkGN6jIM1
5KtZAmgwBeGgYcscFcwxSXTPrMYTiVmXCQBk7ijoeRNLJVmFhL/T+Bqbtfok1DMxqpqLYDqbccgS
l4UxwPUorY7lElPzMNlyxgwTYbRopMBxETr7iDbIeL6WHugUObsP8k6ZIVXCSl84FmXaP0z9ZJ0F
aIks2a7Ovau3ft28zYuDJCfLwcpQut0VYC+qYQktQ32GVzj7/sPYCzL96STfSjEW5Kz1yJUUJQpM
MscFTZNjCR/UwY2NTA8d56abvmEukogKu/YaQUKcJ7gEMsCoMK3p241hrg4JjjxDFrCC5m0Dyhhk
uNfwD3v3uxtJvkfPyFKGNfZAjq9WC0oYySXmcrlqcpgBLLA+kk6jzKH92ilSt/+pdyWkHyeIDAyD
CucRPtwCVuhSTD34UDe+FmZHgzlr+NnirPtwcWH+KRAD/TYyI3d0dMmXQTl9BTW9zB5innE+479P
HXVGltHPZW3QLx4qZci1s56F/OGRkwsXep5SxZDw2icy23dhOwckcR8GqesOy5XHBMQU3BKTKYB1
4qB17dlUnLQH21J++qIqmn7UdwrbQAlJPF3DQvJS7lctjj8YtBG5RY+ju7nK88x/CNvnvDJMKJbl
BO7IL7MRoYF/n4zMHkSN1jXF+6CQpmYCMRF6aG5C7yyQkU9yJ0GU5ZgGqMUAik0OQ3wzz23tdehg
fmBt7v4IFtY7DX2Zyoel/Oplf2GDlYqoHISVn2pbhej3iKVE4UjkNBwc3EbJJgPQleHpo6mJ+HKB
v+juP9MrSF/H6kg5JRqtfZ5x+eHEEVLPPc1TwLs6Ud4csqjetar5CSyMb8JjabQflnyB6rG9NxTR
/Emj7eWUgIAzV761pQgfC/Vd7pmWzGX8LXEWTT32GZUWaKRx7lrXXkI9MasfXnr+rFjBNJjZSy/g
wZy+h9xdOOFjXnFlF8htvK0Ohfit9lRHqifEc7qC4RVuPFsp8hkTxIHJOhRiawQyd5MGqwHOW95g
8mk9GAyA74MdX9ik0xtLFWSTHlJS2Zj7Qth7VU6Gtg/8opognqu8LPZdY4cdyyjjMZyuKmvTCeJh
VtP8iTDq7/o/YmpZwmTT+HACPatVXBmFUqS3kKBr9tm/6CvKx//vHOiR4XS/zDdFYZNYs/qhBB+l
8aNgW4v9dTIyXRlmvSL+PsgzY85591DtoIhCRqsS80McSPu8/CNldc9ysfOy2FunLtxrAkICioo9
QPvxl1ieCGyFEHsxgkhR4/ajlD1Yy3jpNrpHeE0II/Mr7c5invTsHrsCOBT+K5NrDN2DEoqkIrO7
ZeZdTDyzrVlzQ6D/ENrEp/pAyM/IWsFVp1Ocw8+bBNye/y99YwJBHrmLpKaKq3HtG1VcSZfed0pc
KjjEkXKR12FDIwB7hn8CSweq/9nhbj57SVRSU0rlsHqznfadswm/wHqpJmtkQt9mqrxhftCI0GxT
SgEwWwSy68N3dep4anAV2/me1KvJtuLXU2oVmyDNC6r71vMjf+aoym3j5COEkBiftIntytDb8MZW
1vOFZWNYvvbDXXKGDAtmpIkg6s30AYMiwUWwKhSVwRPz/6EIntb/2tFVhz59veagjEhkipA4Fbec
rd8e6tbZ8JYz3tRzvzse3IdL7v9BhjFk3cACDg7fCEtzi9Yd4I0vVPSKiuWJ7zF01zHrgor9Eojc
MFzzkdf1Vu8w7t50VClueZV9vXQZpedmDAVYs0mt4rMRCbLxt8i1DPij9sYaDeQzNuuhectperZd
couaTI+kEnrgGbgPFIlgQxXFp+pW+vfudFiXc+VOF/y0gMLuAA4qCmPUmZ9b70Ro5gHn7S77Dzu+
VJIAX8oWZzxMDsg1ak1ja7xxICD8MNFZMCN6BPQvU240mM4Gnqb5hOwwRotXWwniu1cKSC5gBiLi
Bj+ZWRDgjq4YBKnMhTcammgru8xuvoMXzhB0EGwi2CV/0QwDhz7vCtc/KAPgIO0EKiKYqTtCKHnN
b6Hc/8szLB8z/GXqL/0N5Rna6LDxzDo9TrKyACAvE1EMq5DmLnbrxM85AYEwB+VPGiLIhEgdxG9g
VGcO4LUVyTmhOFzb9jOlNrmwVGbVMQF8wpKJSxkyDWTnCL0oAJfBuzoGLeEZWIqMt9Bp4v3pl3BW
V5NUw+F9gFLUntYTPrCR5uPh5vHhktkVhJhYdEdPfFORfMCdU8HvQs9pkzOA7i5wBM1Qs8wdDN+I
R8ulwJT2AqXWOgB+nt1IDIxO73yHNdEc0vEWsZaOioR7+MoPYMAJRWzvLTCEAEyc+GSO4wDvoLZM
4jLQXX9TWrsvVjRCpWjrV2jvapfgbQimMj2EgCfWoM+eyAcvDcH2G/ZsOx+AZNhea2cRyMKn9ZPC
II4gPP7IztCsDFdebwv0/jDbKpKcS7iOV/zggUcgr4PX2X8OxLB4uf1spfaNgt+Q/fiaE1co7tpo
sV7Domt69nNsnHnCUIxiN5BYeNFr/B6XiZN9XEo+tHcd91qzyeOHy00IwjlMNbY0UhNX8XaT9dy1
2KnL+gcizeI07KWzfcaXTt7IG9+L2i/MdRU2yD25TdErEkOQYtYBpDxORA6gsY3UOmod1YvKKcUh
3aIMNna8wxX5+pJZCkbF3FzUXNkmnywq65yBAujHkfRqVAqXMJkZNPrV0wbaBjpQQl28zt7PQryh
a6PjS4rkXRTBkli1NDJIAO0ui8lOmN3lUQhcG7F+nUOtF1bme7/LcvCqP6X8i3Bw43l7f1AjaRZK
gixHhaCaUYHxiL0o8b5nsbpoQTmyq9TJFJiLfFldpoWPhE6YNrXS5R44B0wjpJVLoRdKB4FIA+HR
Pm5khtFbYSGDGXI70kCcH9KvNtjgw67XGLx3bLdvS4VN+fWJBe73RUfWCL7AaCqGBuV+LU2pkKjF
sIoJyQni/g5I86ZkOXWiVlqjt49SMn6p5AI0DE3V+N4HigNacsFa3PoAZGrjSk7chdU4t3G/SoiD
SPk8qW9hG+QKm4OiVTEs6MoOgTfHA1vNwnpWy2liWwwAmb+KPsXDIxKa7kvrSUjw7Fp0KJx2fdNm
RzAH2KDZmXplfdM215f2l+fjBFHNJ+eLq8ae0PibpTlYQfoJprULME5pC+ZThc7r3IL38FpHwQj7
tcke8cqSFuzR8RDjp+Cdn3kOBaOCE22J0j6vJ/WhV0f2hYwbkZV9UEir/R4I9wf2pxE9kQvAm7cT
MqBeRyy5cJy/zUtDpxCzYseWnyQjcopu7qaM0hHyOFEpfNJbgFxHZzBKHLvzRoyA/xY5lZSyd2J5
DF9VtALxFzndselQheRpjfAfhWeomdH4HkqHE0YzfTJ018nuHSljuBscNZjiQlu+yIASGTyxX3ys
MoZU+jItEMG2yWSZ1K0DkcKJ7Ahghj4H68De3k5hVmqR9/ClQ0joZaDSay62dwA0iuAMGsEhtyzf
7UbzohDPXZjxjvNDck1nTDk6jFxXMPHg3gDnOY37kjZzmCih74AVYAXJHlfiSLscECJAjSRX6uNg
58j+rxqNtNjo3Uk9I0ztmYkiH2yjKhcSUceocNo+eEVWF7RkTw/pSE3cOsk0HQY4Tsx9HFsTr5zc
U9uyqqGsbHaE1EmnSU+dtvVC17STBDVEWfy6OmklLIi/bLSz5VfUMnsxMt5uXvwrKNFu3oTjipIF
YREhbh9pR8cZkrzkCdnikg2EjvyMB2jSKjRkmVZGURKZDFsu6tmtNz/haWZ3EJiO6IDvL+TUUa5l
uQhkUKN85uP6m3XTldjctVTP0EvNvdjAMz5/Mtj/zdD7zKhl7WrKU9G/ZFVMnM9TlbkpX7IzZQc+
xWwcpl6Uy6e4dWSxK0M7LcVeSspvimIvbloHf0ndHfd8vzLNKv6AsS5iL2U8zTZDOMgQSsAK8AWX
kuNYwHGtGe/lVNS8vcT49TsqyHWpgzn776pGX2XgbY2Nb/+v5+yDCT+9MF2TDFG+47YINOOyVQ2f
js8vlFDNno1hOVkK+ozpDIjQRkUViE9QZ28flmUI5cRBU3zvkPXGXLRlW8WxVJ1DCiclJA4X1Fbg
2lZUYZ5v75tp/ymJrp2rOZbnr4BTZ+03nFx7Hb4XtgFOT9Iy+Njslea1j2YxCpLDJZ3siNw4x4M0
utWOQdlEcwAyUlDf6aTXdkdD5LT4sEiiyVL3V3wo/WtSK7oyWFwB1hhPLkCqdaaKs7a6Z8Kd2sjw
3cBdYQCg6PA4CY7Qu8FZDL8ZGDDRZK7ATJtaEabJZlDVO3sHZRBcywAVug6rgHF1KXYdVWJUjlU6
QWfRd0d0e4h9XGv1/IuqpCq82T5i5vjR3yaH5hh8kwaubtgb9HRFqHmQyS3byTFc5xLzZq026Ngk
J1RAfhunhuE/EX/r8HNVFONcLJjIA4uyAEzZCVweP7PPzVxgwNve/noWDqtuxQrn04DoMrCZnDX8
jOrpW5htxx3wLcMN434RWFxAxqynWGu+Ehf4M8qpGO4fLnGYxkirAXcEZvA+9Z9Y0R54zVRsUujr
5yYKULinevEBpfKoRNWpGsy4NYFQRx4aXGwgXvW+XfTnao8Tq5WuNTb47E1hOyxel8g7Wqr1BQoY
Dtsw+muNhqqt9Y0329WLxXTi5ACV93i/ZlOOaeZea4UWVYIKXhFjDjPn1SJzvkQ+DDiOSfPAYeCy
LQlebsDOGkX8a7SMxrY/3WJ/NrGamNKnoYYnj8Ykm0tgdtNiiu1OaBgPxv6bejNq5GDQWcL0CSLP
Deao5u9SkJMQoG1hv8IqcRyd7yEgQmpjMSwq8OmFiKoAxtvHXsJmUvmwgtsEkAeeTzcjMTmROHic
bJGmCzYDJUsAuvIqiRlWUYCe0El4xo0TM86B2cwG0BYTK8h7VWSzEdJDfTBlU8Fu4IJvH6QYVSft
nhgnMrsZaq8ETKw/tLwys1JpIRDi8iPXl5d3FLgqqZOQTZcpcLT1NgIGkBN25vkXqTX+vEReg0b7
NpucxLYYP8rFxwO3fBLxncECpeJGW9wWMRFU1/3s2gcxfipTQEnp34hTCrD5QTwNsl0v0206DNpT
FuQl/q6V9sM6qwHNCGb5MzvvLRp+bm1OctgFyFruW0rkVBbPfE2nxTuo6NJ+SNGty2zxmBDlAQMp
TGUYx85SvaVCA/bxQ3UyiZ3IADHMxcJgaYWyIk9OYTPmVu1NkVhJmadcErB8SqNyZtIW92dwi8tJ
sUlryzgVzC+SdKlZd6MF0whBFUW8+ylL8ii3YhKs3lZ3dvMxPpcoQjoLh/jcGhUfurVsjTn1IUcf
BzFS+yKE8KYlt3fne+m0KKgTlFvmO+AT6BQx1rPKhT3WGOivXil7e+4SqQYkfnKSLd0O5gG1RjMO
VagyQ3gTrok3Ib6v+eEF9hzH+EAuFQr+3YoGTqfBRUrorYO7y0ZJ9dKHbExUd45/d6I8vPUZO9/l
E8bVv8b57CHXvLmAiaPA6/haa26DCGgexHrMgHAjWCq49vEObuPE9fzYU0+v81F9ZhMn+ZkKnzag
JylQ3rY9pnyF5KFth5EGyZhjHqRjJNvboW6yMLPXVXGyq8xP+bkns4avpeFC8oe28H7S5eTjj97e
4YL9mSDWrEGmJwm3roIiaM6ZsZDGVAysVwbIEa6uLGL6DAkg0XRLOZik/JPuWfsDyGh3DaZoy62O
+LhZe43ol6J+bwNy3KNrzO8i5r6MROMQFC9InFZD74dZzZeZLOIbfnU/ApUwSI4JaFIqP9S/oAEm
yy//yKRhJBZ3gmaNP0XaRcfrLYhOWdM42882X/d7jxS7646UPYVnA2mEzLMrABr1IhoJcHmEyVIe
b3Uw1bYZamYVN1N/jCFbZTt0wwBzAR9ZVSbDpDeJzrb2sk3Kt6dIYF2HqGab7R6xmrFz7wBsGXgL
eTyC+UorQnPqPG4wm0zh9JF/pb1onbloqv4296H3570aH6YxETfPbSXypavXGIdJg3LKT2WZP8OM
pIjmFhdSFXhqPm4PKBI3Gw/IOMG6Jmbsr0npKfO07XAnCPbnRIeHx3U8BL7mAwZglOe2eqBpo3wr
SDeF/7L7G2AjKsPT+I6kjyWuJ2RB7oU6Jq3dbNMld4r/Do06eC0x6W8HY6b/rNtUJPcdlOycgKxk
KthvvifOx/+6dw9iSysDUU/1lYZIYsl7rgUVSqARXQfWHi/fZeC9xItRvPDV2n+xGCk5UCnfplM8
y0y8948Yn1VWfZFtDlGfjDKuiddjeAr8APiKjxeKoUfpQf+bcVxnsibtOF0CD1n4ZHC1RJBdySj0
iGKTjVs933RvC8Zm2figNzAvJn04F57jICnaoF6x++sBss3DifSbwifWqHoa0eSSjx1ykYOm0L4f
Mi8x3hTS85gEeVCYp37krwVEYGZ6Qx8yyVn07+SBfN3LhigJ14VGznW143nM8Y+FsNNvJSV2PdVt
eNwpYOj6rYjvNX5Q+VH2Sk5B6guTEywowMoBkL+VlyF4ArMOHQmkU+1o9iWaZ4Srh22NDG4sUsuL
qFVwaOMLg9Crl1IM/9jm1Qm4PavsLZxTB8Ke4thvpjK7awux8v0MYwCM5CoRpyrmsDTOnBEODvZf
0UR3t2b5/dAFLUPznQ5Je6Woe6BRTRSBoM2A6/IzCz9SupGHCswQkFcIPmVwk22Nuqa4a/rSRVYS
W7/2T36PgPo5bKzsijXY2ECNcHn9d+Ud736RYS9KfESvkcKZf4zT6xZylbmSYOdOGYyCEJdNiq7J
RXsfUb8eFd+axMCAd/gy1CsrnSru4H4FBxrkw6OyJK4QPzqB3TErrP0mOptS8fI+cz7jZr3rb4gL
PDHN6qY1kjXDUIr9Fjk9QugMUHFxtIf26DbM39A3KL6euOLK1wwyvXAar59I0lPE3BSQsPec0BsY
5h57b4fAz7NoZNjEYTCTdJ84741AqP+niUpR0HbixoDu/MmN+NJ/7toddBc6c7wCOAs7ZStkIXZo
e190Q53mZFPRGzYkRmIKvY9ixiSyMbqekMtm38bA/u7BsPVS/rFL54UkC66FRggkUAgK4LHccJbF
GagCAAcWyqMhVFNb/nARmlxwuz/DgoTJdVlzAxiKDuy9Fq7VaYP1J0JyWWFO6duXjumLlvjZ+efi
+YJB6uktYZjmD9hNTA8Gb+qX9hEUKOwVehlmxDujnhb2q3jfQyBp31Ljf/ozFu+0MPEA6ZFw7qj0
3ivIlqcxBb9v2+sPjQCaU+d04Th3MyXTmAqckGT9BeIZJz0f+nyLIX/Ms7LWI1FG6g80XjlPut28
8q+vIOkqs22NEgslZVm73sw20waMq8ysqVe5CNHG6zPQeY9PgT8IdZDAnYNf8U0x3m3TuibhG8vA
RpV4zsE/mu3UCiXabv0JrRF6geknPCdVDnHLXW/bbJIeRdAsf7F6mgI0RrCGHFg7RwqhmR+R2jgE
9/O0CqKnhuU7T2hn+q+91hvPZLeirVqYxEmtVeCi1pVDqz61Ldxbrr5t2Mm0OWyWIxaF4Ze4pEnL
d/PgpNZEm9NvDa/dSZ0zZOCkgo//5x4NqBVw/o7UR5PkolU5OjKXO5atULOw+NnIPdwrKd9h0P/S
kSA7nBCFINL7QgfbLkX5QGndx3OnK0NGzwGtqvI3QuJ4PWTFaekOGuBUN5ZwXs34ES8iAKO00z+C
jBJsK/onY6Pgm9ULLolfyNyM3fL4VSntpmyU9CVnN+viY7QtsA6JukmYPG/36SP2/4zeize8UQME
VnS1vA0/wSP9lki+Mra6M7EZtYwZMmkderZp1mP3MdKGJO2v6qvD7diVuJnPaEHmrvf27CYRMooK
8AhrteZUiEyOImbmmqvgf/J0E3rrqMrB1UrYWdsrjW1FykpiyPNLyEypRkdssziGw3okrcOvfd7x
DzT6ecPa4KkWaLugUQSPfzEspormC917xsjhyBwgj+1FJXQsiaDB5Vwcr3GSNtPrCXIbS+EaACpt
PPXQwWPznFu4z6gkn+qOydBEbNDcoRSus2lKC7k1nI6wCeMK+AM/6ethC59SbO/PAK8R3Po0Q8Cm
jJQxFEdZ4y9eZILF+5puyjUV1eXmMBFPlfSANRP0LdyOI3eAHV8KObbdELB1sncHXvhk48fTXWzR
ZxSs9p+h+6i/s9YVtFYJtrFjZOvaX/aEv7gecgpfxhqkPtQH6Wvykcf1kT3YaKVifLwcmMEl5pWe
US3cjI/ozYMrYWVfc0RwFPgTQ7xb2QgY5o0z0WtAGBMTSC6tl1vn5KMhLupjRIwex7WYJO5MAWhH
flfZU3xZnTQdUlEHilWBgLvT2iI5Hm5YjRcFjCeQTEHJQBty3tTN613Dl+0shqfzM54eifhMzKG3
hWiEE0LfinGn6xs/XRQOeZXgpq0/FqHKUvAoKiQOZC01wNSJ/Oztg4B+CKiRZecp6BeXokBYNFXG
fpRJmxNf9XBTqE6wnzggGllFngZfUG53LT7sgVbB2j+F0uDzWXDLm4WdST5RdZqHh91vMW71CdkH
vp7Yazpf70F58wzo8s6Ci22j0qfophPOqxPbEBmtvAzgtsZ9VEU0rNbJrs9dagvBhmUfAqYmiL8G
zV63SVAWELk8WTlH6iPw6cSBmpsG5X9ONqs3UuNxHD/NMt7YpQr3n4xq7XyGq/Kfcyanb/JREZoK
b84fBp5007J0hJHHP61p/KPTxpFcVTLVtyAELjMUP/ylBIJO2FSb0xeNUa6MmEzaK4eUDEhDCqDz
YeUZoV9DZGmChSVSIhPfXiNoDlbT3OxiSuc5WHA4/i9R7BvcrP2vCJr5crN8cdfgAAn9lQDxQ8h5
NJXHoCBtstrzrcYI+2IxlRskqJBZGXxbSiWfPB50h3b6x2OmvHF67ntLpiMfY8NX7xo1huPveik/
blnCoi/Ri4SxI3Le1890UIvyR1KekM7+mXAMp6ApVaEJGAvPM5fBcnHAOIq4WvfeVzhyl9of1Q3b
FNjqEw/gdy09PnG33VUBkxA0a911XaFqf6u0Zc8LChTVo4q6Rj6yYWFJnQuYGrMCXyUagaPH23hR
x0ocmGDQThHtWhDcQOb2ZVODqggV+g54xE3xyrkwewdiXlaa4Yq3oPh7jB87M8/e0HIt9kE3VMOe
cV3OTNnPLX8Oc6Sf7qc+7+V5V8/yG2g3YNCXM8fyOCURHt3dXRZUEgMxZ9I95xyan2VCGLhgKLpe
Q71QiRxvk+fiHuDXPSER8nfMk1EDP3UKoIH4/KHxCYM0nkTX6b+zbSDhJlcJNzCRa8S7isTTXBeT
0WodeTfP0qNNTxoJwOm0Kwcl1ibsQoYwnp4vvmt7ryTvlvr7FPTbB8cuh+txmrTgjqOptG35pz3V
FGUx3OrJdKz3xHAzOM/PegCtfeooXCF7IqM7+k5BS1SsmQvuzY/kEnWOkwSxvKJFs/RIUvDmh8Em
zCtFVIYCy5FMWhcko/25pazeAql46+Tgd6STntpHGmwYDcXAx9+YQLF+z8svkI8AWUb52flOvkcU
lGw4JI5nmA1WwOATeRatNXVCkdBegAhq6Ikn8/vnS4v/+YDdcOibuVnPJ2AyFlzbfUs5HOhz+HUu
AS5t1ua3Bd3Nj65SE8SMH0fc+jnInbO+wi5kvvlTcfzPMalWcLPMrKt4pUQ8yiDHxx35Au+RVmda
GAXagFNfZZ2SARu7NouaboP+HJ0EYoE9ZWye77ZYgkw8iGuV5xGyazJ4QqCvirL0faObAnTFhWpD
VRIXLVWmNZ2KdEG5vwMxQKLxFX8Toiku3bleh53y5Pluy49iKEH/7wBQEdFDv4dJ1HtcyJQVDgIj
8ZM+s2fgyXr9v2Zxx4bL/8/21lgm++zqdZMIs73/9LsSUyT3y2F27RB91Rhg7CYROFft6eT6gG8V
byVuvuuJJ9h3BIB39D/tBM2tlEC2HSqzsaalbeL5KzmoAf5UtjOIHd2XzN3F1Seq6UHZ9SnyzzPJ
aUKpgeLhv4bYP8tSV6hXWD///Qk+6NoAdHNK4XjkRcoyGc4WcZWTjUzw3IgcNvKTgqs7/K27i/G1
IUnoTBCLSVwkm8H1ZH2mDT6T0Y2doAgLHUmcy2aqvNxoBzLYykFepBEjdjBljz/w7kVcmykqIljY
SPB29JJHciBEkYHEZTIuKCUYdnDtFFYOBxPpTvxu+4aMLVPn4/c2d9Q4X+IvEZIBKxlNLG2iNb5V
fZjGw6Omdohh1PXRuRL5IfgyYgcPbtoY8t6/YokHcoJfMPvoXHvTUMlFNvTXSmZUZWyQT74fS5Rs
uaYtVfhcQ6/zlNwF4/hPQ03EaLV/FYmMJu0tZ7jznc20fMhvmylMuZsQ4BK8mfYLLuKAh9QzDkFs
pj3Y+IDMiCSbOTJie3XqX0AGgec8/8pvam1pTD2N8TWkW81rRw3d8wKIigPMxNyuz9TO+WeAk3gb
Rjjr6uAumrpDtMa5HUCTXyQFgTq4mekKj/Y1mBkAIU6xj83UdnyCiLCAMKfUxW7FnAFmUCTfzLlm
eQS/usvblUjnr/XrIfQlpmFEAc0BOhyQtyyVHPBfCwHypKYo/QJ8lyZdN6ecvHZJKb1Btn6MPCtf
xZwC9LKApOpGLZNRSVfVHnHt4xCh1J8Fo7y04e8Jz3yuBQMMkcetEtI8q6tHCsaxaSQBx+JFaGKL
Ol7DufCFG5DVsddP6vfkv0BOwkZox+W1QTGS86J18Pdrb6wPQmF62SO07+r24v4BzQ1nj2wauyJ3
SskrfABOXhaiTsiGTy6irGbX35xZUt8/FU658YGUwL9PyTk6SkMjLO8kWV3w996nFQLBvfaF5peP
hs3gGx/8PFneAUxG6T7xL5/RMjKzvxdOf5p9+EtavwJpKFjInGuW64Cq3+sjQKjY3+TYR06bSldk
rlxGdmfr6DhVmJR3xEZu516SyTlcqvsVMhEYUbi0w6X3k/DO7kj8KEELiB+MNHSuxovLUG4MjiVK
UhTb9UPhio1P3PbHrBMYRlaotwe1ANYyT5BGBRVDn8kGaUMUqX3E6FmZw9WEEQRgfgjoSkYuTE2K
QLWzYqWGLTfTh9E13yNsiV3G5nMKSmveE8K8L0PxzUWaqLpoBlADvb9hZulqs+o5GF7/IwQPzk7k
e7NOszRC8CYk7toecv5GBysbjsOh9YhqwwrhXG3izGxdONtYA14JWwmw27mUpR3YH8jNDcy2wzyY
3RQryhKPbrd3uCLIFQi/aDNNKoIbBnB6q19WT1S7OcKWdo9E0GiRq8k9G5pHNrUUpGfxWdGBi93r
YT/t+w0Xt7h9yKTS1v5NzDntvtckJG3IRukuRsbuHkteJ/RA13nUFUCEBi45dzV0AI23u3FdNQzm
wTwx/RYfb5xql8HhPpFxhBzncuWFiXxlKgCxZOmpGFtho9M7XpFRHqSs1smk9PTNXX4+GGMLFy1M
obZix2GIcPUlGAw2jgCe3TCPiWhw5uIhnfyFs06aYn5S4zHgyjOMJLCzDB7N/fPBY+psiYEOj0aB
b5IzTKHP76OndY+fZizWFi+zLE/SVEQZ+bgC779xZr6v3v1roXJ/5wtP4IvT+7wQ6jKum8T9wycD
2O1OGmxJewEWAQhqigA6cd/qccie0l8c4G2AsRlhekV+L3pX4AIzPCb0pCxAlNG9eOF0NDISb0dW
BWc5APZUgVZgna0yRPiQnZcdpRpunbCwIGE9Y3WjGMa5iKYFs3s04WqNYitH5/eNwTeS2RD5DMIm
hzSZzP6Bx8D4SdqIvtbxeU2TDrdsJanzHNkTKtEUDgtt4HwJ5vKIJrAjb1w4Ufx+x4PxMHtrKk1z
VuCSieCefnMKaMq1fGuflwZYlsP1enCXKuJYa+FVx06ZCLgdrFZ9HVA1AHgWLkhBWiHpXUv/Dgdy
Q8wdk2PqJFXg2etoYgHG78gQj5y8HyyCPqpNeHBO3JItMXoemsawYSq+Or9h+Ws7F2nLkM3nuyAd
hlfHRHsvWykTqX0t9nLmTDxQjvyQLWyKcLR1r8vf5T+Yw3rgFTmiUQmyQDcPnvr4vHNCyeKkWsDr
NALUv7ToVtMB9q1XVa9pR4A4iaCprIPVG5w9txBTJvbLuVCXd1tPbElQYTn/GRWBhEJ1OLaBU2UW
/AfdaVsP1Ox3bEwVOdvLFytEX5HEtlEcMSuE5JTCGhvjMHtWor8Ap7aW5/1R7YRgDRHlikywEvNU
sAHJydmQD1aXkbi/3KOBuSA8a0zk0o2LTYIrLEGcIKP4fp+uurAcYj84jlpDxWZww1Nvp3DQbmAL
gtb9ck2M42zMCMxjMHs10r1+F39zAM2ZEin/JrEWs9sIr+L+VROELffuIr4RN5yGdTdaJ/VGehbI
A9r44nSj6WycvyJkMpUiKM1o66UshQFLzFhry7yONOwjKxAAG9NF3U7P02iGLCAa9+jKylf5lQea
4o3tVdb3K9iGm/WJI4llqxoHZv0i3jWTzEhniOlp54+tJEer9YrCldUpP2kY2ARPwNMNVK76V260
HizE2JtpWe8Eu6JEeHJIUeJeWJOcECP0uDm2xxrc0IUJYLb3YdEvK3aHtZ70Aml+c6tq/NsV9oTs
LOf9VwO4D8CrKdYSANB4u+Ur9WCU9rpOV1iAHGDcK/zpKgqg2KwYtMNlUAupH1r0pWdpeDN5teV3
KmLmaJdSQ3i581WwMJZbZte0N7pxt2dNQqtWRT0v/nDiDkyENj+dZz0FmJRe9ouQKoDFIJlswIRg
g5tJ3dl4HIIAKMaAg9KWRzRD19OUB+AiARqYXHCBKh5KVEj0oqiqRZygn8S8YR5pmyO4n9pfr6AS
lOjSxn04HMAf42Az9svfg7piN8CswPk+ICEG2LOnmI5GF00aq4vUaSJ4r5M/nzETMHziEd3qeqaN
Trm/D4ASj2ddvfW25ULFBqIEYhGX3MKe5SUqqAhJZmAAiqg0co0oK2UdlGn92b3jn3/veBnLAVSR
wRYAxts/Hw41+kUhpxHgHF90/G6+7vm89E3Jz3omcRkogjQXLTh3LgDdcUriDG25tVadcfysI4Uf
O6N1vh5rIuoMdKYc94Od2QjXPIza4O4fzy8xoE/olGeAd52vrDt5g4MXVdJ3LkLHJ4CiMJbkZcD9
gjdKKIPqmnDo8ZwhtrlKPVliYb0XfDkYsn7V+naW2jGTpPUEbBHIi1urhCX2tjWs/sB1A66VkPHC
YoiMWEISy4gSqL1rHzraDRdX1Rllk586h5cHk2jfuDz5InoQuZHb1+fkgjVarf3Te7lghdHHYkR1
HLHCy2DlOiqaRSRME6qbUTQiDdmL07LcrDghenKFdz1kJlzXtEH+1RS6b8/SfDf+P5mDAVqwDnW8
eMSd9ew68I+wyWNuEet1ZRAqRn15oFesbdpWfyj1F/9YO46Bi/1qJTz/cV1o8Kneo+Opc3RLyhOw
u0uQfWMwLpOiFEpWihLAo5DlU2dMMU7RBXxuwGuA767CfDTmPNFDq4fDdklmtrVnoESM6zkEzm64
R8Vb7UEgSVMaqQ/c5DP4Y+PX4C25eiQBZ8oX/dVG2yVgiDX2l88UwWN6EanFAKiro/jddXVSZ3w3
IF8a3dutpEBLg68yN7sBu0g4Z6ARRc5J3ULnvuVf7m/Z8s/IpkJPSBsvpKP9P5DWL7Z+OSa7wrND
UrWtTq1VBwfwrHPhu3mJAk2syPMsIKoBRdnJHryrAXX/6gs6blMdXAEW6w1UpxarXS/E6+oRDQ7d
Spf+DpDI9i565DkDu4TiIJr/2xlwB2jB/FG0urFm1iFmxTjopNkPUh9pqqvVvwSjdN9gULrUYKR8
YR05kRJH2saXU2an7o3TfZ4gtszkI271GKGPRaOrpJyXlsHAhGVQ5XHxEZLI0OCFT5pBpwWFJTlS
4zPz1D37EQ18kXQTYSlo8wxx5blJ8H7fzi+o611YDecZzYgWZcnN+u90bk7W5+Nt919+k1rMoE0Z
Z/z1Zo9X885m26AqeDV3bwDOadkNVNMSJZ/0SipEH8Y5RgGkRPFC0Y53ovTGoNsr4jCExHDhMbGy
liBhWT0yty+15kSLFJxm0pWBZzqPh5KgxerpZUmc8Iwd1ef/LLk+DgdBzp/FMCDZ33aBGTL+hH/s
xfGgv4u0ddHR06TsQ9N9gFR4iibpMN45vB+hKkr3r2CdbuS6eVMRvn7uy0fim9bFUFVg5QiBkm9H
x34cPE/FGUhqnenZ93fu8Sjea/BG0CDKf6/Dt/qle4V7tY7RrX2aMGU73C/RL86J5HJl0GTrnBCv
B3dqfonVu5Mx0hr1fn/9kse6ncEoLuu6KHFj2KMyhuG6FcYFemZU1ACA6ZZzaO/MHl0LsABJSt3S
0atxhT9JNSjNN8x8GZVWWnEVeYd5lUprz/u1sLLNTQ3pgyLIcKuCyc49hTjQ5AUH34cHGWHGFBbI
4PZS0OMjXPuhCcA368xZDjuOyW5EFn9m7yeVeXVjaz/5PB9GeKAvphCfkIE5QyyeW1UlKiqMHB1u
JTbW+f0R8aQth6cFQLnYTWoD2wVvUEqWRvH7CRyM3UrR+Gug2Oo2s4wb21qjxA0eQXEDnetLsxbK
FCs45gOzTbKpmxsgIztsOleZ4K+DFJ5tFbQromhMhBjCWH3whsM4aXZnLYs56PLGSB90u2T22GpF
BCw4CuuhEEHMfbQeKmrLfv02gsWGDbJrdUAkcIeod3tw9IBzQF1bTU7agiKn6diPSPFvoSj+mbwL
OMwxtKd0Lhzttht8npQJqsCmLiEQe1B3Y6kwAhd/UWoDz2Cro9brFlpazkM7/waZrEpfe8xNVd/p
ZE5z4Zf/KWLHsmCa92Ic2qbhXAvmApctfWF1FMrZi7neLqgRWwA9+NsigA+KOiBPFqbS338h7SOz
ArbiULvIPxezApVpBJRev4YFX5wOlp2p8/otQWg427QeK+FU8Qi09evUK82CcLha3gXXjbQX5J3R
U7FDiFLBtb70t39p7HHfa9OQRg4kxE5gMu33ARxyiAT5NypUgvvW/4n+R5yhmWFFIPx2hiOUqUT2
6M8oHDWuaZhVnIsP88RhU/XgRgGeRc2SApk99+1IFdCcxWJJuJuwXefWeA+1Zdq5HA8w7oAQewN0
jPGXXzcedy7KDPhBgjs9f66IIKaQkoPLXlCICnEllOixiorQaN7m/QRJVV3WdSn/yE4xjNn3fE6D
2eSNDwvTsV6F7LY29yLpS8dhfOmOvyoCrFJzHRKIVxyW1GnlQ67qWmZcTQIbrzljeoZnMf40j7eH
bi79qJqMmURTJg3a7bbwtv5SVpYyurR6b25qirnMbwdVWlWb/d4YcrBARUH8tYYCSN3rM8Q++9zb
LPd7ygAlQZRCjgGPCxZnYbtmHNMgaMa32nywmIPWSNybkMIC6CP4R2hlbvhhZbLJSqo8i3o6X8JS
6q2eFZg5ZCkJnXg0w9SE6VTn+jRwSwvLN7aTLtLbOt+hWXX2Gx6a/vflen7bTqbDIu0aLmgAJQ7J
gzUI8xK/Zx4+GgFCilyzOsNm+rRXw1uRaNJH5ynrmDOfZBMWeViFJuv3Cz/ZSmkPYDR/u19X2FYD
1Yg772HYjNQoAwYvUYGbV4/dPu7dp2PKvaZeV2VVzD09yeX9y/ZLXOQEeBFX/swOyyh9ah+9EpXy
qEnv9074BtH/iUXT8qYhwYgZ9EQ9ogZte0IS7h+m1Lq3hcOo5Sr/+/0u9VhWmmAILF/EujBdZSur
2hvBrMuXSTUk+vVcmc0svS7G+Gmb1AvDQY/ZaJvuKRTaIylp+LAAkYyElCf74fc90ApSmChlM1p0
VFmsfZL1r7GZqGTQlOJpLzYT7YnezWfw382WKQIAPMdcEyvKnoSN+SSkBGLSY23+97gcKc0Xp1ZW
0o8ckawN5R8/FZWStonjohaboxYZtqU3313cSjpuVrAUyNXdYYx98W4YN+rcn2JyhZ3UOzGCcdQh
V2KVKJ3XyogSrvzmbK+eZXhqHqCvdZhmmswolTRsWdXDMg+6FNr4cwUWI/ORk/US4GnSM+ZY2y5e
TMBwc/Q1fth8FE25eJHlZtuCdFTvMaTT3eKlB3tQvipZ59HJhc/4CZLNk2bRX0iwbp5+a5lETh0v
oBjQZ4Q3Wq7MInDsmB181i4L8Jxm36mXgqOfbaF4VDpmKTWNibsiCE3nHxLg0/0Ecx9k8J/idleL
q7knhyPs5ZjafHlGneZbYT3QcOtsRnI/zNG2OQVsOk5T8cUSt+uif2K6XOVF/eMMGtchWACux7Sp
cABYEyyL/bWJ3hxa2sENzwYGE034/zbL0OHhRMCfRFpojeLsf62h78Kv1jHaWd7s/S7La9q3ppZ9
zbzHlLp/lHkaggfHMtiRRbs10/Zbf5J4gL8H10cWMrooxsnFCvNaAfPCeP+OiTk5gdSGqr4c0EBw
xgOVhlEosf6m4LiYwxi5hNrVVFE1s1sUJq9zYKzzq0gdDjmuaAkXjLLuHrSEqWVU5GOmbCTwI0dX
R3IfnPvi2hrAF5Ku2cyevf4RSV/7TrC8cf6FsT9bcAgoCDmiuq0RQEdOhSLrioIDzPnQ+/ZSmKgh
37qiPlB2owrajUmxAXEf0GyH5FrL5J+1Y0pMSDRHgtXaCqK3WY3EEe1wiLDLIdRYjk8RkGTkpsCB
WoqEIa6nN3lu20EfWPIy/0Bqb9RPSvv/XLjZiaFh4CuMlMxLeByJp5v+fA9xsEdB4o00Gdzr+tZh
C/gXwDIsytSaUdLgheh/b6gxRazRVWJpNcjrGYhrq3O+Pofwc2vi0hzrtlGgfw9Zh+guubGFFT3n
6HZXBIxW6eEqdLC1SFgh+Axw09i41341taZppG9NgTPtc39pnWbcuNxmHhZjEbHuRvoWGj4ADW3+
zosvfTUO66vv/8v4GVHm56o5UqMy61LTQmfW+T2C/1c2HTmXOpBfQEkrKcyxyq4JF+xPWv9wacIn
Z90hKSb3QhYzSpFxJ2Lat3O5wPJudRUDZWXgo1BloRKWUyVzYKDHJC8lHg+WMWscmKHXbKYmAzkb
lGfTrIKSwaT/N4JtTe7ZZYA1kz9I0fdKsgcWWZfmaSuTCaONWBl8jOU+zKRSTZ2Zg/B/Mr94oXRW
4FRPhOnuY9WoWPIfzuKuGWI0+I3nZnHJk+6+L/s6BDvmgMSDctakamKWrFfB/NTLlLV1+/y6kXY+
oSMxn3TAlEGReXW8ehGQ0S2UX5wmSKg1X0/wXY9ztdQ9HrIRhPOSTjiILHdcJNFSDMJZlBigkC+3
K3bheMRS4RsSiDM21OPGQZHuWmlq6huo73k1SyTdXyxIwf9SgmSnazm4ApzgpnVBD0RZ9HRO42QG
l+IaqJc78OiQgrfu7fHDLuPOrlD0kfZMPzkGiqU2fnvgIMvzkJbel5zo2ByjmeXUezVDpWxCxHaw
ndnYEbhxu2Ry1RttLDlspG5rpQOC+Za90JAY5XrNJ61obpfcVpbYdESh3oPcYlNDTeQztnwEJh8z
lLuJr9za7pDlOAeYjyoX43Hqj/8w4VycTueXDa2Scrt31Q5EieG/+np6qqLG0eSnZiRoDgZgg548
NW7G0BMrruSzw8gPGcqlQKiAJyqc9lOb4EB975zWuDgqL9PeOt9atlbhYmaotkcsOv7kNkCV/HVZ
MqvQXtbyGF0/HxsIQXUrR1h+3cZ/DdYDo+TuGEbqnjbBDy8ter8KMEkRtDXH533PlWNWmYFclLMX
mOkV8lMjH3o4bRKC1/lCSdrHCYb1hg1/b6Rygt8JsaE4ZwWPd5JSfCCrh4g0J50yIHtg1I01fV7h
c6Mes9eSD1wRtdCAb8jtyzfHWP47VUq1UgvfZFFxh1Qi3Rq1VLf1wP4McfkxcLI91cjFxX5EvfsV
ZBQexMyex38cIjIpUrd3vEgnSQ/TSbxpb+Vwf58g1OGuQVJnRgayxzD3JsqCVYucSQ66uBmSYy/W
cZ+tlmvnNKmlTGpM04eoXWvs5MBdKRWKqpRBYGSuNTsAgZtwsl8I8Dunt47KqXfiDIYwAAamm/zF
ekO7n/a6gvaRru6ZCa+OLG6XP40hklgmEFnRflDc6xEXc0sEXd8M2WC73dsHG57A+WxaXsFJaZjs
SCl99qP7rlALFOuqjA8ikBSrbX2Z6PGzvn+xeZ2ZktE6va820DX/28WOas1sk/d4RgWpo76jz7al
J80TlPWud6J486tdDnaZcT86IOAtJg1Yf2NrlhxHC5UL3VTL4basL+lCrp1A+vhNWkjSs50utkWf
H/qSeKh5FhpEGsgUsxtt0uO/R1l4TO/hYmRd7CPkfpzzGm489KSx+mM13s2iumo5P0SrKsYpKU38
GfchKa7Mxs2lQ1RQgtzOdasXgecVmDyQzllqkSly63RwhJgkrTjCB3PIlwldgFqz3ZOp2QqXRgBx
V/xFcMdL86zeVfPKJAqZWibTaJjsv4PubVhdqm75jB2HPieTnTxOVvzBY1wb1TERM+hE+8rWPkXQ
/MHJ2Sb/X7/TITikwY2SQyGTXX0yjGRCAq0XIPRlHLNmAN6NX1CJwtQXcBHoZaCR4G5tRge2yo14
6IhRGuLsBhZy1jE4F+Ph72DHf1cxG+qc4CWW3tZwTF2UKJHopL4uw9nr/C15JQJ6dhlbUdiM8Zyh
wZPt8AUwWosO1UcdGRXeL0I80e9deBOm+VVZYzeaIUcZ0KzN+kqW6E6F21mgFJoile92s41w/R40
8lj/QsfbiCKywiN1Hgc59pFJMESloeilOkGHSpsz346wMDPoUr9A5HHvkp3kDYOi0OgWzerJF3oy
eovwcxebtpoQo7sFOu0AacsdguMLUE54uq9CcPo2YTkYEC/eQ7ohC7WyR1/lVyYulmT3o3sustqy
CVUzZzKv1uqD0nynEuzAt2BouzqTNqrFXXGAyAXvobJ7O3APJgJZoBGLqKq17uPLaD5jAfAysZsc
giCnie7zvyLHlNNgvCxfQgnKw/WVJN5sr/b8jx7Ohzajhp/uHPl7YQwPkQge74yZkjjEFRVlM/SP
0RN+3a3C7k0Fws8+oK5Q/UITkpuOBz4V1+9zM4NaOM8FrQQSp/9Zwja9juA0cBLgehckUvK/+4Ij
X3RHCrXNqo6eXkqSKvBYYBnGeVy+KvKGGLJHIIcQO6CBGJVLX82m2cxV+6cnX4BVf6eBGZJiTTNs
HJIiKcDx+Cy5blvTFW2Fu0O0iStVxcQXVn17fK0fDeUM/Cfo1DAASpHMdQiHQLvq8X7/F9wHOmbb
R/yZaFgM76LUuPR8EMxeW42Qy2tKIjVsm5u2vMoW4JxA+Xg++nLRqi0VROcL7HghsMSb+5kHqDZK
PvpWZ6hi0Mu5VQv0GNozcqlZpjHONZbj76oH7fHaE+1Nn1KwYOCto0CVNw8T0Yi3iS6HQknN8Nqd
u4nezarT1MSaJXoxwAOfx0YOt+VsQtdCJMn8HXaBNfVLjhAwIGsbBOAULqoE5gAjYM1auedBiDRY
foM597pwWa0dg+6q0gwlC/A3wtnhg04xw7GxzPBOd174AboxkCEnjBOM1P28pecLSFMCzNjhlPtY
s5PhakfJc+iu9ihw2K1aBjkU0fV0JOEUHxISHdwbTQq81ce+xiMhoyYoSRokfwtjxE9GA6dJJiEx
OHdMagrSFkOur59ZFry1NGA0972M8Z0yEFL3JEiarM2TGRUOvQUcffC3LC+o2+aPhqJFL8t9E1iW
lHdRjjJ2GHYq6el1wiEIetQnefEruc0Row/nIRQ7Z+xqdNy7cqchUbsAxYxTC2+CNsFLW1VvUxaS
tQPnPFgKIFqCC8Srr0E+j59LlI6+qtiyhzw/Z7ssUkS/mitJLQtFtLZ/BoKpwZ+BWbl7gHfW1PiT
LsUDT3kVjq/OJutT+UiQw6QtfL/oZb4Lk5BUO8ziXlAyPqSUXLAtPyz50ky7lwDAZ4iSG6IP/mS3
WHQLnl8JybfsyORh/TXNVGWclOJEGVRUUNo6WDCYKu4/hdnE4T9CrwKBVol9Njscpt3plijV1zfQ
tsS689yRd9pqnQ8Cq4/GxO7Z6Ubi0rklqj6FU6dpvI5jiWjbq1oHwqZu0jFQl7JDTSRuZYb4edk4
nRTB/TqMu1RNhU/jxmBkOget2ytqWUZkj1lSE1/AXmtJ69Lf2ueuePLANEXy+DvCh1Q/fqjMiB5D
VCGzgifK7ICm1ZPsAKXrYlPi3Pr+lxsaVB+Y8zJWTuw2P4dHF/wjOMmQZOfhi18FOyurY8gJaa5K
+dyi6ZmS+FsLuAHsDMJiPZMevjKwSj+xnFeRfZx1dLhtghzWhRPPU2thqwG4PMHkFzb9eoZznIwA
6GdTQTGXKN4r6FiIL2uGl7vjYhwnDusFyefXHRlec1PvZtR+FvOcdeB10OCDzG+cZUkInkblI2sj
c0FmzrpHzxyCBrlapIdsnTwd1MhAZL08InctsCl2TC+rukKtRODcE5YxkdyhJ3XrDuBAp8qqm8R2
+H22pUjw6prx5+ynWoDNgblCp+gRcXtY0/XKnWps5tfWnEphH3WsoS2dpQOcdIWkLDslmZ5vghkp
fCeqYtBP6ksT2/J3bMSDyDrwABRsOw/ikNuPO4cDUlAhHx/11MRgA9dyer3UnO0DfLgSlf3Siima
SIkhSRxlfWTFS4kltK9Kvuqd0N1nklC65qcqf8Cr+R0Q6jjOWyALP7PcU2Zjrzmieilv3KEck5k8
OX6HiEk2HWZXpyArzMTCO2++0YX81UTIyy/eC0NmluuaeYY2v3tSoouE9462U8lL/+mxXyPscwiR
qfGooefJiseVFkP+TX3tfLTiIPlQ0TMW+ZG4InvqA+Plmn8mgcPpycV3FUxvRptlClfTJNdZnccY
OjictlfkhpWCelwqLcE133V2VJ41bTwU5DVmhJjMwN+JrTCDF0njjyH++zDYN/8N0+9lfCaoqtfO
aseQuUkSomJoEL4JO1NLH5nmDeZ3Uu3vZZPivjar1r0H65kbkiN8aE0lU1OaGxjSzjGP3reL/3vy
u1vUpobLGRP12xZhUVPmZ059k5vjqWqTTotiqAAGOvkaIV2LZCYOmg/3MNxj++07tXV3J7nurZKx
TwXVwrOdJmwl4BpbBJUVuJUVNNa5bGr4KCbEQtQLRysfnPcSfEWSybkBniwK1/E6dqy/iUx6UzvQ
Yr5jUo9mIdotkVZ1Xqp2FF5Kwx8zRLJVS60PEBJ6k7fBML5wtmXAOKddCtZTkBVFj5/l6PNPsTEt
r8o+Z6LbTRMRl2fvXf1lzYM8XiguXyOUmWvWn9kmFExkP2ddOz5rVearuMALpCescu5QdyUWzBxQ
1587Q5NBNmAjx+VvF1sIu7Fkls4tJt0NLyDZsD/ihYvmRn2fKduDh9sa+FMZI8kMJ0AVWwZ+bnwO
YzI1eYGDEKE4peQiV1A/XU4+IUd7p25Arg2mSM+jNq+qEtIzyG4XlrRdQ/Uk8v6SZ2G1H7Ut33T1
aYWTvs3RXmwICUrlLEDz6nIlFqWguM3aIqViO0jLJBjbKbfZ/M0K1C/5zp5YDI636nwCVMRrC16m
ZBZ1ut3DxJrVXDoSeGQAwPp4r/soXOOYKAsNy7uuFkQEWkcD/LXWfo/jE8P0m3HcEgB/Zjn/iX6r
3B1F6j2kMdBueq0mbdc+j6ec3j0k2tF7+Tcg+oPgKNflHhkyZrnbNFcnVuF9A4U8MllzaHioRJcc
hW65bGi+NyZiFvIv5Omqt+H2tFm+cJgrTJy2cRX15tW3/e/sO+6zfrrVDgRAlc0j9/7l5jUAZBg3
448DyqPYDbaQS27RSj7Hku+/wJ/AdC16P5y9iZd5+mV3ZVgfFBDfUOM7vmf5JUX/MN5EQgn30iRg
Ng4WIP+R5sj1CqEFBlM6bU1v28ZjZNa94/f1gx9eWocmCq8jsCOKx6VyHzeTkaKiCkKoZJU9g9ip
COJOXnReLuL9rTGSfFPTy4JqeJSkzZh5RXeBpCtnxnMNvnJZF1gfyUBzUyuSruQwzQs7vYZNmO6m
ve9ihzde3PoDB49FqpvdapT9gTFZZbiJ76BTgmND3N2yUUHIxkPBV3EwV8nj1DB4vNXxnrlxY8tV
e6AJUA/5HNE9CAVkm29vugsjAsAMUMkDuQKdc7WQZKlUAZ7QgGFfr93pLCwfl79nbjujIKDoXiIc
ufniMi0Y//u4dInKNykFh7QqhROQVQEgwArrY6beMhYa+Zs7US18r6KG16MVzIUjUcVzEW7SUfQJ
Sbtp9ooefah9jSMG1LhgYDZNcQJF2le8nmNGZdCE5ZzioidCFz1gR57fu/6lLs0xo/aT6KaIXdOb
JSf7V5FubmewjcanOJtdztK9pt14gxviihNslnPT1nIYysVfl4uCzmn7i1oWMX09Oo2ccAJCxS5h
E7Tw7t5k1XMmNKjPq4ADxIAz21b32qpvJq+kL/YktqPMa5wyOejf69pC5Ibl8lcVSL/cdEHL5b9L
f1iuFTtdqIenjCSlwAORU21DXz46JGUowQFEzFqUSNCTwYV1k5iLczX3mC2OKQzQwQg8hfj3DmQF
5NmxyyBT/YldXHkukX+lscA/Lmt8t25oV0VZGD5FCpIiQ480JhKcuHNT6C4aMr8oOO6Vm3W/lcCz
V49IeqQGdsIOqZV576monSzxvimmhpeRDiOKDvDTExj2S1PUbKkWsooQfnJlwDDyKJFKCnnxAjsS
11i/nU1OAXUgsLWIx756BGywp282qhS6aEpVZz4oU1fSkuE7QurWBOlMyze6D5FCCwWPAP0bGS3F
CqNEP0s43Z1Buq7lJ9yudRtavjBiJ7jKzb8Gpt4ch7h+hsG3wJNorHEOkvSkyB5yREC16zaez/O/
DfLB5Wf4XfaB+VQsy0njd//HeZ6e838bVg+dqRJUdtG6cEG4KAizOupHNxT/9XgL0/JBCthGRVy3
P95IPpShbUnr2DlpcgHYv4rh5l9IBC93hGCPTtk9nDQ36eWfRyqJdEt42/+H1JkrQvBJSoO99y90
T6yeSXkL4soEN0M7dg8aiNXcZThNRHEV1KIYDDYjrxUb2yw587A2U4pNYd6YcxJMsAeaq8ixsz5K
+6AST6VUKTfOA2E5YPVsYvQ+XbcATdIIBX8a6fXm7t4D6Xd950ZEisHqNgpq9QMur3QiMGYdgjJ8
ttnGiEnOD9oPQtFqY+2W+x9PgxIeAjQI4KdaPWtKZ3uI5VYZgIL4mqrW2qKIUafbAPCGzBOTAeXv
8vAIWe1U/T9jZ9h6m5J/LOxbSQqPSqnM5v6y6Jikq9XlcYE+mOQq5HpQMKdj8rYCtg2eSyOx55Oz
NTuXqb6hQVCprhtdnhy3HLOa3HuP+QkVeK7igVr4VDtWUcjGg4NJK4UY41dlHOQ/KsGQ4mcv4p4h
wrjs8sqPNIAw+9g7AJI8hRWJCtf8OqLZ/oGDbo1M8X5NtrrMBzVrKEO5nG8A90jMPTf8qOHHR/p3
fBj0uOgXpy/h2bDndLG7NG3J4CGfaVhvipLL+kzocZ6X5fKTY7VZlswBhhH3cLC/4OE5fL5ZIocH
fp8HH6VGg6SB1yZAXdg9eVlQP94Oub8tLwqsm324BsgHtWb8uh6EGj1kfnYU7S+unUE6h+c049I3
u32RxERS0qQwdXx9maOZyA+U2nVGqH+JPBnRs5hJ7i3cg4tRknjaqlT2T2xSSmgJniKO1QC3kpgQ
wXhRtgD+JzpJwL0BUJBnD4BXz47cqG8WkNQ7ortn1mn6RRp+FZqUaffNzup30+ECxb4J5jNaU46I
a7Nx91M2A7AwGbWAdouOXXXWWFSWBJSZyzq+eOCItS7yV5SlSVDQ6CmDepV4vge0z2yvzYQ9Vn9d
82Qp/u/oq0pz3zFe+L3N/vgAIFB/u/1NKYXn+whRjYDAmKCdjeMD/8x5t9lDiY1vt9x9OgUCRJXc
7HuwAuf7BOW1QOTHICimLXNjLbGkMs9I80X5e7ZM0BLh3P7lpOqvhTNTzeLW09DITsZLd7AxKIkx
TQtHlJ4DCaMvpslawktcXJERzdFrA6GmyKaEvkuIfh/aWuNgiqg79Gkawu7mzLLdka0RVgRuXC/a
VynomBo2X+M/jV8n77nnUEJ4p6sv6HgY58U2j6blmpiaJb+O+biHcJyOMrgFjLB0o2u5GRw4BIzX
Vs3h03X06ZkUA5oRBsq51c0espl03JD/STqn53wzftUH9PS7aokDSqY71Np6aZnXxOmXhMThBnws
Ho4FiJpHc2GMWPjhzqvQ5BtiMbQOlfb589t7AuG6NM7juW9SCsj1JsCqxuDoKWnJaFuzBGo6hCTw
Yus3Wl7kokAegvX2qcqH5St/z1z515qYlENfoGvHJAzeVil4hMtBh77zhicrFIpjQGpxXcEf19J+
JZR9wTNaF0WPKRw5hBPstIzF5/sGpNdeLf6xppjCPYomrPyZv7Pf0D/MbRwyjZvP/14fn+5or8x1
F7Y3613ILz2HDgDgi5f+3peW0At2E3eYdr4rmY7W3S7GWWAx1fwaMtFfK2zmSJiH/PNETQTxblo1
kHbP0Dl5nkaVMpRcoUlcswt/7htmeyGk1ueewAg+i5efJA1V5xceQ1wrBG9J3n93lXZeeM+azAow
6TF06875vleP0HhdVa6oexez3fzWSPSBCQ9oGQ3r3JW0hjVo8LBNByTzJs70b5Zenvv07Xi0pzfP
/pLPlSLcYB5p54eLNO8dbfeizf/MpGTN0CXV4V4zK/HIgDKvoj9BtW94krc8nvKHztYywGFroXz0
XQQMXokpcGJ0HTBk54DcGJJDAIJ+7Ec/rNrWmr9EbthMxr8vYbsvqPtY0yb4dI9mk6fN3aYz1l90
QcDHw/pFYYknv2cRc5ErG59o3/Sl27b1vTqB4wFoNaUfSXotDX9329npMNtQiwkq119wdYyIz4Kw
oUNQn0T3bo1SgZqn8Ai8yro1sTdwphJEBa8QiCEb9Epvqlb2bo1pvoyuEBMDBvZlzWS3uCVVWsKA
fvFsoDtHeYRE++aGbQZL/FlPPf9gWbqAkx+mWNxFSYRo7h0DfoLFKsM9JcRBVRIceN7LCubnSBKg
/POgESfvEQhorcwDlzmS0JN0SBxoRT3KqhGbPKudS/Izdsc2lncaFLIIo+1cxu51YePrpA4ntN2Z
aAOU1S/0eCB4xeNzAtupuweHsEdJNSoB0LAmc/LoDjX/KxxmflPGk8b1fJ5MyctCWaZ/toFR3GG5
rRBQhVTUUBXaRPVVxdvYtwYbf4WVUDJzG+IBJk83mEyzBxdBqQBiBnU3Sa0RH0JmMVxMdXQfWC2t
MhHgP2fIvMjBJpPgirCehCcEXkPCLbxBeC4dAouz0sKsLzIFW68QHVecxLc/xEarl3H/CFYZNotm
WQuGY/8ZAgixJrRx3u0z5stVslcd0/27J51kSrWIFHeMqurrXFK1ymXflDCPcEay2BoIsyPg4DHu
Inf5+nqbQ9JQpzz4zBcE9oh4gIbOkut4dUABSJYnEaWL0OSdfFXMRwfeBiImrAg9+1ZiXBU1H2X6
NMb959gPqxYWJlnZDDSmPEryfklZzTE0idyskXqIGJ5rlP0+85/5nA2UTBHALhNZiJ5WCSqkF8j5
tb9L8g8M78WxLy7AkMtd2rttpTgXpsu3CoIXv9bspWgo2ka0Rm9lpVVk0fJzdjkDgRRyl1+Iz7f0
ItvJ4IoiBK6McrmonBzEnW9VHaZTzgzAaZFcJp4qriQksn97h2xO+9JbHXGngXeoRldd/im+xJbM
Th2WCQEzb5U0Tj4kbhD3WjKK1X8rGsb7JGtw6j0IOI4qjFsSZThUijTqPAe1F9T1LgGX2Z8KK0pY
RXk7L7YaONBQcVpXDafxpMYMAGMXpewsQlVXaFePLtZmj4qhcd7pv1vSQHCeYaRI/AVttXK/gORt
2igVcwBQ3/J4TMIjvB8pFasl82Iro7Zbz7r7/RxM8MD3pooR/CfwVxXoHfciUO66pwPtaPJOMeUP
YkQtDMwPbkAdtgm+ZzeQSryguVAeHJ2yt91Jr0KnHxuyAd9AGXHLH5T5oR38xeDeoAFSnU9KftsJ
p/WSyCwdeCLqQJj5jD7H/LTLMJyDdBsDwnM0aoPHX5LZww+ICGHGbFEONQXQllAyPBpM34M0brmD
l5yHrKy4902di1QISU+ec82M2wzdGG4Xi1myXMykbdGFPSW59KhtpEt4cyWF4yOhXgUtYwGYlQyA
GT1kF33pUI0R+2v4SLQd47c90G9sCvtUMXyA/BmIr/Df7/lYi1EM02l4C819PkVaFuFdoW3K0AwU
tYSviXJfEBKA5nIEoi9p14fWuIvXBGRrGjdSA4BXwp8GgcoJOyD5mIUYfVUqmgYqFOPsMmt12odv
yVBs0Y7SrQv6FTjjgukTkC6t+bOhr3EpmaoHaUyp6DwBOn6O1Mp1cF1xT/hNjOEE/DAdJyOkwuGY
FuAGKBqaqt31o9Wmvq1iAMVk7m0AT8V9rjrEEOkW7L6jwrS1vURqaz94iGLzC4LiO6hmuG8fcp5f
dgCsMf1YQYo7hztiH1N7xdMGGiH8QSPGmfwN9Nx0g8sBWgmYqgXgVojz+n+mMm74gAeTJig40PSB
I2ueOrdtlnVYp0V7tG05IGeMLAdXEQxaAIBFb7uPXkonpTiOs57vAN4XS3eCyj2PJvF81ZM55p0F
PMK4yuyugrZjM72RWJizIoXzAbKwTRqq2CNHmRdOYJfzMKG5/Z6Hrxtz7MlvuhFQ4JWteRO3yW6W
xXZi/n2SOgqu8Pfv+z0tP76BodXxfDSV/ORXZ7Vv3SAdCvF5s4/qmuehTZBPBWHphHmHWuav+FFf
XwHjydgfGdAcG2xYSSgyzMVyyLy+rnPT22YB2YyHfreFQE8ju/sXAf16eiGE9LvrjU4PKweA9pRm
NFU1USFafAGNVH6U4RhQZCxWN3ULleCpz7mmPz0MTE6cxtpj7UMspuUxyTMlCuacFHR9C6VjKzNx
B5Jl26sWbUxxdLu9Keqg35YxaFSA6mCfBPhH4VzXi3V9VchLtW4x2OlQ0uxpq6je47vmH2np8lsV
yJXfmJESS0C9qFhUiaZr2LrgQPmB36S5nx6pIn6Ve9A5yOGt+/vomPHjdLI8iBBDtfKlUy4cfxXH
ephNY+CgRxAsGoHMoea7m1i+wEWOk3NYgJ7AmrgEhnSUp9EvD5Oh4Gki7GusUUOSLyFMLWzcoPrh
A8wRTxxq/370YdJYXzUqesAwkNfp+9eeRUU7nELq448NpYBal/HR6Sw6sXUhyu1gENkSg4MQLAHO
pi0nZMVfseL3bILzC22WVSJ1nAja/gX0kggDCQ3ifCqISBQGiRmbPynTJZTw+UjQeqzmUBehsIsY
xpOgqktaJ3vrjes4SjwGPhYNBSWPpVNyQrno0QpaYOF+2UvmOj5vfRJY71VY3AI+VIq349AHJ43r
wmO/A1/+buOQzw1yysk+SdMhG1a78ummx3jqjwEIxEJJ14FJUME8oWEL9sUG2TSFGb+1sm92/qod
VNVduH2JK2z4Mb2DRDpRtECymOoFCVGIo9sJDMi76dd/g+JXzqyL5QLkVgIXmKanvwk/qKaFJg33
r/Faf1NWmTM8YHaAb2MGW90meyPuIboKaIId/hIpRT5F2o7bgubRLnNI/b9ilL/5ZUU94ljSsG7t
LWCkzOqLd/tokO/QpitxHsgGtNW1ShNqLfxXHwzSI3rnamhK5H/RFutkL5lhQ/uEH2uWusoopzLY
m9Lr8bPgi7vVvn51qvXlMtXMzZURU0W99bXZL+KFppw6NJ0Oqt4mvYiI4PVoi6QUvJslIzHtPmK1
R355BZiCHNgNLZ34vRpcGX4rNxCP3YuA2IqTXNal1D/SUnsuwa/kKptCP4n0Y8YKIXnNImdJCqJn
HIe5Lt93VZPKtoiXe81q2ljIz8b0ojk8jPaDCbIwo5gWg0PtQ+Sd93Z6tsKzwcWCabzGqYc3+xJg
REUwdCKdqpyj73foBNaDp7RHdIloCA5V1ljK4Aw+6HWkVcalo/asmTHiHFRpZ8QQT8vZpy/IwDCi
iG3v4OKUAexRWW268s4wU3Qul81rxS5+MqMe2lZ9AjkDB1WO1359m2NeB7p7I6Pz2WoyM+J3zASJ
YvCLUyBsqNDhXKJCLyFaWLmanoqX5Gd/n+0pI9W7KO5+ZCCZGVSninTuWm16e+KIBAtMUsbfOGxR
fYShlAELtF/DAszx+UoKwJ6t73IYjg1nMfzJo8mtAcrWBFGgvkyG0pMIHUoz9AoOxZJWQ/rsJ008
v29DWSS4Dzihw3p2aysi32yyRwfDOx/YiasperlJOyFQ0pyOyD3iBSrQ8bVXFYhK2bbLNYNR3es2
7RY91DXmxYL3eZ9uRjqxsugfpDlWdztCTXtfE6npyumgaWqAYJl68lfdDDKZ+O4VJwqc9THPyyp6
ZcNHj4Dy7UryIzO3WQOebrPHY2p/uiegtzk2jTiX9PWyYgHBhQwR6cU8ZdghMaLrCHKAJ7ZfdVZz
H07WlOfB35y1ts7KIdWUg5ganMkxebOV2X2G0Eft1Km0BSc8c4Q6A0rGnaJUzjK9wcUi2luofocI
EqSKjWxOX728i5qQOmHGaR32bjI6yW1S2UFCHwYgBJriRl9lk/pMHbEQGiWMQACEBWMbWK5Aw0sf
kNlNiDWV4t8JJkc0LFzWilNaKIXpSU2ZMcbAGZe6Kj04mmaDfeu9lmzeZe4lt7x/8+suTPJDManK
izYiyA7oWpnPiZmXoE2k2Ds6SbAGslpuowPfk/DF5m9WsWHRNvkE1IcD+R1GQffzsPdiT4EjF0J1
xkeuMPEJy20sg+i2hdsP3IL2EqNrD0cNI6+hT8LjT0N+tXwhlm1SQxebVTZDj4tFIrtAlD+rD+af
Zeomm0oNqdKS7YSHKrZbUg76R/LUKaerdbB+ryklgb3ym+g8Tdp1CYsCZoTwjw+h6jzh3I2mSTGi
ZEu9WU9dM9/H15PULKlcPruhtvZSYzIk1lb3/EN9V9P2Zm7WA1MzaJAcyVp9xNMGRH477mxTa+cv
nrZbbZ71y4P9JO20bYV8JFZmdCBP98qOdkJ3N9sreQUn5994A9A4fuYyrGGoRoL4qApk8Ux/RS4x
uir023KvtEdWbTCFqmXgNJQ3ElTO8upTqf6wYW+/EI0xBIyw/S6ZQ/K6M2RhOf3rpKggMMpWN/4Z
nGZCe6BScNqzEp628h4ncA4PuGZzr6AtfaQI/+pJydeVGOMMl6jrCgsLcA2CGokpmA8kFKvWcupy
KNpRlMyGNRjAEUi3ZzuLeseom4Ke/0Z9nBwPdzQ5i6yQ5uQ3eY8lgTuLEd/t+077f0Rm6Zu6zI+/
UmuCvPrhYNSeaUT1iriKXuL96FRHxup90sbuzZSAvrDOkKG8b8kUWUb5Q1kaCLtX2ZtrTr2NphpF
rrNDe9UiyOE0j2CfLBr5hOayzNz0gwOwXkR4VimbRGvOJBhptwqEKxqfXFoxHmGnG+Sqi4TTn2Uk
tu4EYPs+TlfwEBGOHIYnKilnawuoxOJFiIoJf47e2XMWSvzw647u5yptMn1OEapZO5KiNLh2iH/K
l9tzcBOBfNbPZiHJJSaY5SrA4xI6MiOcpRHkmRKTME2JDg64SM65THE7TD0reR+waG0VkKcwtKMk
kCVRS3NbHb0vSIfu3XsmWLEp1h8h7eU2SoZaNiiRr1gGh1m29sBlO3Hqln8LT3nrVpuIQCStBoym
cWr4K3BrYdVb9wyY8V8RBieO6zfJYwHi3QdaFmzzzlqS2xgCwOwYXavlTz90Og+P3Z7+QvGz0Gdz
nlafq4tCx5pSdmLglxIrnpJTugf6ldsDFNhQCm5Juk+5cRLmeZAwpCzMGNuJUFNH+zA0bwnTsvDq
Op7s6DR9MfYnLzJY0I/clsfqC9Xo4obNZT/ajSwnqzeHRHYdy77BK6MUFG3ohM74OpHuinzM9mfz
9OS+V0ZdIcxrTwzuI8UbEIL+nQRLsjFcHF0iHvH2f9Im9wFD7jX4Nkf0ulDahwB+z1x8Ain5DDvx
bTtBBqRiU2JB/W9ck1m7bL6WaYar8A4fk5D9VbVTWOPIpjx/v5dFwNorUKOLB1Wor16WQ+YwGBcd
jmQk32dSd/p3z6L/mczBEogMuHtbEZwMy7AVvDbBnzPEMl+875QjiDZs3sp6mSm6VEkWcsnR+H+y
FWO8NlAvK29KszHXBcuJ+TQq+72H3qQHJJkPRwcy8C0WMmy0+8Mx1SQuSzraEZmpp6VLGurKW74j
9qulMvsf9L9HPpXFaHnMgv1/Ig1kygF5fsjshCRRv8D9VDpcC1ddxCfJcS7ErVFJ+46Yd5S/vAnq
SmzBFla8JXW8cXjBz6cELeVnlHx3pc/sZokTuxgM91ubPDM9OYA2M9WEercfL5huM07FDI22TT9K
o3xrJKkVT5H7TXR8EiTC/2G+dFPpA9Je0JvI0OL6zORe0P/NB9WCEU2wz62yqrJHhRQQMyatCdTh
qXvt23XTkDCPjG9yCoQph+WdFIBycc/Xsf6BzxkVB9eYgrMfG9Pe/qsCHp/79zCej5NXJO4RGOt6
M3cf/SAzBMU1eh183qtoqRmfuP5T98W+0+8mzEFvPGJhJFTAzOUH/RF1o1cM1hSRxdUTJSL3KuAT
SYd78y0fP+lUQxJQXVDGBXRyI8ogb9WDG2+2teBl/2FnPmDwuZIWYW/d90BYYK4Dnz/gIe03Swbp
33Ef4us4W4S8Qts9Ormpn3peN/0UC4+kMmiAzgHxQXZYrS/LslPfu1gDEipA8fHP1FN8+dTWWkpu
783wAF/fFcmQhU4kUf/26SDr/QTR8FfzeRC9suCBgDKggeQ/sTKGbUjG+KeLcskuNvFvoSHHWQE1
rgXtixJU6n7TAftp2kyWd17IIJ4b7qUPUEgJf4v5hbF51nYJ50Umss+murw2C1sEnyP9kOYOdVfU
OmbyqANdqGdu2td12VRaQUs+KWx5CYjft976U6oMixQbpXWkboBwk+tKoFSfb5iLKnXWubbjqmau
Gy6d+BktEj8yjyF4boehTvH16aXvTVe5Uoiquj9Vu53GQhOHA1dhUV/Gc6QN/NVA7KDyzV26LDOM
mjWGILW44u5Rt16FbpBpHE4c6bzAddj61ooHkWCqHHio6v0FQUL68PLKJ9X6DM0wpNByfwqOS4ws
5quQu9XjGf8vqwYGD6jml01N6S3ucrhJfxlpc0mB3oaXLh9QkqQULaYbH6XF1JCg0cpdVYK72W5c
ZyJrFeD90ci4KbWRJsyD2j81jUoJ94dWPhbe3touUgZGFGif0Kato2fe8nMwCBivIUKg7H/3cFGu
iy7Dl6D9N4mUR26nIwbiXgcst7a3Ud28Bf+f4P5WQ4g+i7XqixBK0ahxNWghzarieijduKs5S7Q1
zpxGNasqpj9kM3zHSxXnx1xbwZnooxrTasf5t6YRljv45cs2yzEzXSkpIy7hvVC7jaNfL95KIqu6
JKjqmbB8Fr0w+TfilG+X2SrbHGN8yybok8waD2ZBxyoakN1j9MHrooWWqU87nmRe8fNxiExDLG8v
0ZMzQYVIukIbZz8tQ4LVv0nOOUqkuvCm/7P1i7VAlQewghrPqcnnihL/ohTn5v+NrDotQT+qdI/W
7VEZprqhTWae41aGLnLip3AhSPndlm8F++dJ8w5OIrghygQdFEMmXlgmTOk1fPTS6ih68i1ZU5gB
fVNbvj8KyXzlveonF+i4DnK9u+M0k4aosZSqzj186FtVHAwFy7dfuaXR7yw95wdbUw6Q/liDoMyn
zAX3T0Y4yVn4lHqr/TMAgQ7gZJUSOywavyae0TsCLYj1CRLmP4Bi685mA0vsJCRClJjpV62ga6vY
S/w9aC+4LikKMLX+kv5NOU9mHJTtcCaQ0Kj4C01toqVv1959nZoYVt3iTe3rM6+TsnuhI4yXzNQ4
WBzd8vBwmNfmuNni7S1/+4l9atoId9oiT68c4qWcf3Y7Cq/xfdE/qWqtTMU/da20u1jJYdPw0Dnx
/WAJ169fpBHXCC6iQ+imjaYhulxb4+jhjKS7kW6WAUFQ1/8UNUJ0nXoJu7SpcjhJgAPYieBRh1yD
gL0SloE3cVvw1ynynf2Vg6L3Fn8YDD6cHenE82095idEM2bhYVi+NvEdW895XUO2+EGRtokCQ5G2
o5aECJvUej9tB8NYSn100+ddQd3y4hAtgli0qaEe9Q7PNUICsUNSOcYKo1KaMegNMirF0D4DRCWd
m/BESotddz2LZdzvEknbrOgrwWu1uwY8sVPZ9dWUnq9PSKfV4ndAr1jGnJ5vJbgbJ8qCLf7c1QDH
FcSPg160zzrdpSd7qxl0qyQhcbMhSQjFust5O1JdGBWt+YRcKtNU0neTMlbonjJMOVvgNsgSHH2R
2kHlPXRF1Xx3zNTWWMe2Cy2INOsPOsjBR4sGk1e22BduQQKsFLksHZj5opMPPFeRJjy5FEjUQCO7
bJ3Sn4xy+jeJN3nZWGlNsKPphtYoEKZOwRHn2G7Y2F4VgIQ5Zb4xbVXXjjp3vumSokv8Zmt5cieC
lHR+uqFYTmHvNbJhp4aR0Yzbxkqti6+3Tz22GFoZpZPrcinyEws8invizC2GUz2hvf1v38ZiP0g3
y/HQmGCffWLbZ3/7Ajwk08XmDFQ0Z5fZseZjvBPparu01ifXAhc2zXBmVve5A30cePpwxeNxnPi/
WsaTTqQZb92rMA+DV6i6TVCRL4t8ttDlPMDWnJZpY0QjDOWd+lpvlemM6fCtiCmTnCha4jH8GJN5
Du/7GY6AV5VeIpWzzQmFzFNr9O/ObvGUSYvO0WpR/7Mh8GDtc+TDEMrbsfXIfo3CrxV7KAh8q46Y
ZE7nw0CkLJfv3Imldz1Pm/Y9lalETXwZS0o7K4J9RKtIzllnu1z114AYjXhu2Y94JFmuYrL8ewks
BAB7p1/NQsUTYoc81GsfownKu5gnOYo3kaROnzWBoJFOLLyYRHZYQxlWj7JUVPKm0Eu38tvFUCfB
MDPCtb6EFDRYX+w2qHP9dFWYx0hnj3E5TGRRH9Bz8NBS5D53O4kz/Oq7ov0GD+sLqv9eIq+WcJ87
Ab59oQsUUrpx/M7S1ItwIjYHAHpTp9Cw+fae2HDyQrt4lzi9CMnOXeTexhweBgGmbofjE3sOwKDN
iZ9oda0DAQyg0L/4DQjxNG7+4YxbJQe1cRyGbE5ar+VVhmXbQw4A3YncByEcq6vkZjPgibkOq9tl
aOch7gjkhnXcutU5BbSLRiYHBQh+n0xfMBqOKkftOXyfinruFwkBryrt0fJHwDPjMAm+wP1whcf5
XhW9ND3Oa7uXLDSjGFqoYr0DBXmnMEp9i8xa6aGoj9oumAdwnWQraInPSXH+ZGtPK4tZ1lEED9I1
SIqG0nNovneGAoLWmfJHqe4u9yCx8EYC1WBJRXh8cmvn8YntSDLuIqxQ3mF0eZW3KHlxNpOFU+6V
RY1str2ze6tSxXB6IoRdN9DzA5l+bANBX2ugNpvYC3zy+qzY19pRNrSBzAsVUYRVG5RDvSxPerVI
ZJ85z+TQcK0pqgW/pP95ZAdGAgu3lXTR1A++ydHQ4P1ym7wZf3hCQYozjd8r/3omZs3lWRIa/aK6
yaylyUxmLrGYwnA0plWypqICi1+3gZkG8R4KgHn9jXqKgHyL+stqvNW2YBmy/qzR1/zrXOkVCzfp
MSny3C6pMEP2qksGHcimmkYFPTZJQEh83WSHEThLDWIMe6m8NhQkf2uQPttuuo7JuIeRI63gpgCZ
/nSuTfZLOyhtY7aysHF3IaG2y5EbFuAcLL3kXBpXmT7VyU5O1R6MG3WgRjNPxDMfXvBo0+6lWFa3
ou8ocZQl7fAVbnBO+uhpdKtIeVHdHTtbZpHt2VmKN7Ll0nbvsReO4pdE/CIJ7XXpaDQ+NnVFaH0V
lwKjvtvo0Mmk3C5Z9SzJwQS4XA1gScl42B3OTOfE6oad8N/LOpTxX3hohfFa3dgMl1oVmAwJNSUu
T8L/Y1hlE3wNmhS+K3bjQ1oJjwFEdNOPAGRm4o/hlnoM4r9ajKhnAJlp2h8cVUoNC9WfQiCwMdQy
XbKoM6xDWao8iqppNWDYpFDm9FRafQTWr7BIcfCQJaP348BZHBfaJA13Zg6w6AoOxGp7wiqNrTSW
pe1d6JP/F8AS94VsTPMmPbLrdiHPl1IuNLFV9mL/tCnRM07Saon70rR+ulYSq+SaKdMHEB0K0Ki9
LsOaKvtUKkfBFtXyRElB73oXZgUTUuxCql933Xak6HzmzoEhWb6Ghfi1SEqiweuFnrN9YwzZ/VXt
10L6foTcxvPXsVtmWLfuzReUwIsm5SBZUwy7t30s3OWeJz/nLhV0/r2k/oU0YF68Al8Xyl/Pv2Ah
qwFM0paE/av1jujAreatpYULxshu2tsQF9Z5MkPb2dRHyCJ1RIuw+Ab/T0CLq3c3PWYlxQHSGh0O
ALun+7t/do8aVlkCDsfOt54a2M8lcpop1eljjDM7RPzyYfCplHxcovhVi3yw4mycxYbME8m+b9/Z
9K9VRp5auMjrciVmY1YzO618lZjcb0M9IgremDVl3Sh/YGQMHVx6KIoJYFLW1lU5nJHZpnaR84Sa
P+eSnqeVxiMRsmYawMkD2K8vNFSEBRlfs5Jt3iSv0s2vkIi2dEZpu0Aq1lGYx0EaXvrKfaWE5keF
/zyrx7JyvTGZedi4v/nPTA01++2M0DjwD9l2NZjS48a8JTSk+Fxf+ujEnf2iunMn6+M62zEMFlEm
JCczQ5UnJnL7m0ZssjN9dbs1102t6YnAKM1Y6DCpzJzauEC5eqVV24Rjev1zZ1PCqEr0ILJ0CdUs
gOqY+HqTgE6GDgqKxran+4gh9eMRr0PK3sHC2Qx8kWJ5jUqXD1/+BhYEnSa9Da7YXRKkkCa6Pyix
/Na+kGz3CXCkbNZeb0EqrOV4mvzymdJ8fQABNsO7Jv7IU0AiefX1LiWQQ25zN0YnZXoPi6LpJ2rn
ah6b54hI2EslYpjaApjarB9qoQJrRyM+Sk1LuXLelrcMr0vwoTPm4m+WaJcUgINvfPtm9caiIaeW
ESuxJCFM6Y3v6sXXd52XFLyJ4/uZWXnlF+MRzrnf2aKD+tY2Hdq7pLl8VVVmJshBMfHDpqDClnjS
DQTmeCYI415n6J+BxJiVHMyBEmKp+QPOEVITwwjpw4G81Ki9HpbFGh9bbP243GGJDttosne2TnSO
UFuun58UK/Hb0jOegMWKnfHxgqIIA/z/mO7xPYTaU8O4r/6SLyPaIYlZ4Rgoj/VMLSmy1T1K3LEe
4r0pbQ6ROYDrBAIFGwmjYffkd/CeI0NyxHJrgXDSXqngcbxqotmVhzfmJmvJOJ953cJIoI84tFWT
tJOtcvddXRrVD+hBMKGlb/XViHa8vX/1X0AQoaHrtGXN3zOinXN+/n3P5fBffv/JSKvBLv2f5bAz
51L6cRZCVAMiCdxA63+dUReNIHqTpm6yuNHroqGy/gXZmqDcqCqrMgfdOSDYBPe3hZJJsdUZWENi
a70UX51RfjDJ3ADNbD6S/byNBXNNvSaxXv8pzyjbObl2kGXccC+dxrg/asY92Lf5mOyRX+g/icLn
XMKqBvZSA4XkuM9nuHJmtlwnFACd75OnvfqiE0Hy1ONRpTNAwNyhu2QSvbVTpTWef2t64iY1SbO7
1YkwHiEteBbAWMJjVZJm8pn0mmYB02dZx+NAkwNSS3HG3BXWENqcikRk46igwoFj5eIY4fddHGM7
k1GWxKamXRgjpnsgkfaFlR0NSVkpeo+egC7H5lCAW0992ptFpdSnXhfx591Ex+kbN7ZhVxMUf4ob
kYN097PiHwPUZ9OpHP01gVS1bpaplyV2TPO/OSZXHNwfplZ26XmIGWnD48YEK2jy0DGbYdbjtPk3
x/vl2+pukGW/BR+0dgN9+y4KFpzZL6DCj2O0ZcV1060DHDfldeaO9v83yqfsMcifrkgXflNLD9jn
CYkIpWgJQvV9zK8d4s+Aiohs86VDX2b2UIcILFoYikujmiFZ5/JJitHBLMw2cItcRKlZl2AbtPun
K0SCcHNjOLtaSgnqCYr6qSoGH4rq/HhCJf0ax0Q4Is/g1pTQ92EccVGJCDT3H7S4BQWSYgGV/hWJ
tHEGLlnpUtbxyGZa6tqOwu11QL64CvGzuDPH4Rd1IWL+l41t+QdkA8pixA+uomBLYzIf0gr84rrq
2wIDPo1PsYwDeC+XEuXVHIV6NmzQh9sEc5mMiuuR36nyTJGEx2cqiYmUWFtzNco6H5I6pihG9WBG
m1+DBgznwsorVvmTry65c2smNfdHEm6Yle/2e/PvQe2GyNeLleuo6pLa0r9PVWkEVUxNop7ZO8rE
zmviPEqkhY+kap7Wstf/A49YPVuy3QmUQTRJkC8jBrwzSmqZYEz/+jMNJSET1N73EeivoiHjgyym
QUXmErsouh6zd+dZc/N10cWHOOshv5//ux9hH0uqxn++j0w4PTA6Wu/lCl6AHNSDJDtvTEUyyWM8
bbbcQu59wymMg6/DIN+fr8EVcqa2/MZcLJ+7c6nFZmzmbdVZFgeRq6p042WGZQoQw2ufxy4a2lib
r2ZCquO6qMf9tejFcfENO7dn1+ijziSOQkYM9gkXrWO1LV0XnY3TSsXGJhOnGHQehuEkNdzLs1E1
cE9tSgzH3K2LapWQ9yF5yWkqKGeAOsg5m0rdQqKk3WmaaVnqoUoirtFSZVIAmz49MGWqGreXCedn
Zp/Aaiswf9TpWQrPaFhCyXfsV493TM+fF7Q3/H19OjMhVsZ/J0IaTfU3zP0douat24So8uewsmSX
4nlPzc8lz7rSBfXYYQiSfGQ3FTegflqdPpA/rX4ZT7U+KzMm/OOqSFXi1h05kDYh5+7X0yS6Z1qV
Miw5AUQyTNhboHVQJ1z85H/E7K52CAAZvpQG5HRmyTA/buaoYLib14LWD/Rk6BizG0WHAc0TsCbd
Dno50F8+WtXG+vadFixdICQPfGLAEYSG93efP1InXHG4YTgYvm9FSr19A3GtGvlCYM3jcsVSaRF2
gp2pmMrmBD2zhzljvEBg2qmldxE1bPCIdHIOou65ChD8i9cTEIZ5HyHJ4Mxs44oN7OB5XgayI0PT
T/OGirJURiFTMMTTrCZmVFz/GzlZxvr0+APj7md3v8jImr6VHcewpJw06rT1CPaS3EozGc8Vze8w
+mhnyjMmTb3M4tBsk2aUPtJ2NMNFHqka3Stva6QDgIEiJm1s2zffP1dX9RECVQopEycfsGbwtYHg
KA/n8LCGtvbMoIvbHQ1MZcp3y6paCQGa5sVJioFsuU2mTxqD31w3WF7AdyZoMNwj1GhLZdAARrZ6
gDyxv/dGsxNTxl+CBMfi2PMhH4LSvA/MoAIxBRxBvVoQoEp1fKscoDV3bkmIbC5wxP5HXWKMmaUP
mP0A5FWlXVLyOGrC7kyiOJMDU+ns30wECmyOIm0+yMbwwDJuNnpAoBplzlbUhNc6qfTgrixhHFh/
yR5UVPJw/LRNueSiyvG/xsf4EYqK5fgFqnCytbI+0kdur8nRDwUBJAV4cjoJEMUBkq9/UGHvwfGK
NsWHkTk6TTGP+FZ2rV9dgIHKdV/cO+4p6fEPwbDvU/iqJ6Oy8OyiQ/7a4NK7zCNGrnPbxYQYCnmE
PRwtptb7cCFm6MIZQILriLzAhkCnNgE5TeRFGwcewFdl/vdIPjwgP4Lmg7SRm3z55+sBJYqyHgRB
qXEgtU9riW60yvsG8Rnx6/HXfnZCkvRLo+rDeuYTmyweAWQwjaznyYCsA4dQ2stZmgg5bvmcQNjq
hg4BkjzhBCNuY2ydr+LjuVIPZJyCnKKHm5HM40sgMfNweOwAu6TGKSLLRRDdpVo9CBEpYLXs9M5V
bd9Is75mOgFjqkRBcBLvhxjQ7+AvKsQ6NBFWHcVrSusffYXOK96cbU262PJ5sz8tMyCqcEQGiQym
faHfS97VnyGMkFtIg48fm3xwgcyqssyYBkVqWndssDM1D2FCLol2KGh7vOQuu943PrYifWveN3yj
aPsZbMuJ3Qd9SgbwAYRY9t5LTZQ8Il5AXsrF5EbIgbNLEgVY/k5mVrtPsHKzJqQz2mlLQXzGJG+6
KXbt0z4+qbdMaKlI5U+3EMn6HC5sWtu+M7kjO90+gB/oLqS4Cf6o/rGpIXc6fHNcBHBurCi6uSGg
nSP2osdMrItkp0W6kGAte+H/ysXGhEdnHkg/EPOxWQ1JEqBU/MDQbzSDQSlrbY4fJ8orEY9yV7Zf
sPoSrV896WvUbrE3n3dnpvqrISV5zTjENgVKNtdnEhMuj1uMz7N1JOgX+yACJ3hlISMM8zyXs0yJ
sy7tMPDd7Pv9OxKK85qXJBsrvngQR9XiMLHoV86uHs68TBuvJNxQIFixX+K3+hb9S9/p65DzpEJm
WRHxpY91FZEnQWVkYScHVdrYZ1bmxiYWEb93+UtYOAkRAUwTKCNWUSm2/FO/g4O+PQhgVI71fPgF
NEqCztCZxK02uc4I6PqkyTRYFI1wDhfvglANexnl8l0KYn64+1LI25tBd7PAETqtcDNDqMbjD9O5
Vmm8krR3coDlfWHhOd+nZgf0PVsRm/EIQSxWhiAOLvAmuZjdJ+TmiX+3nDYZD10zxJwsumPXZ0bD
ijC5ibvLCoaSaTj802ry90M93avlB7LkgSojLtElFPK5FvqUydp4/Nk7/pOygoFxM390z1+sMQMT
Wfztbao+4qyFXP6tfdWFr2xoh01tLUz+yk0BV6FxixP0nwfkVsvsfxWcV+hWd43HGLUt5cWzjsTf
bYJyeV3mesz4Q2ZAUpDbuTbx/jLfD2RpsZC9b6HZplwXu3PTBlS4f85COcxcToBV7FyMgRpN9ab2
DIpxZmRtPpPBNWdfHWB02fVIipCHerIY7UOaYgKkeXcuWYfUN9NcKygYvY9O6zlCO1YwbhxowwR0
FNCd8uGI5BwhLPgLgXxvJUPwaebb7PPYLu/Nkw4cP8HtSuQ8v0R648Bbe7kMrwnBpcOqJZHmHLWn
Q004p8ycbFEp3qDhz9Lk2bJ8ZPRSWDO0w4yG2Zg3pkxu8MucmS8LAeCxDUZPnWbTaTk0FjKPxVdG
L4obW0sXUhG+Bw0/yPtLipJHuOFi0p9VjmZgMBLHdCsjfyW08x3de029KfEwKuvvHJBi7LAnhtOM
SSENQjobsXF/3Rk5hA5lmL4GAMv/shLNgwuVDL2+GFQA4DHojSW0mTuP8WWmyHITSSvUlIfzAQvz
nBOmrQa4OQJErROXCz9hR35yi4M6pDBPVC5T+HTEqIHeRcnQIaZ837L8HlM2oIpEKmJgMf2q9cfA
w0bZ/R/A3vCtHeOKmiuwZBrOgFqEJfLYGGFxoo1SCULhwt2qX3xsVOr7o3m/ouGobGr+tPmOnZhR
o5jlCaLYUSEUw6yVoxiV1gAXCMLRiSfI9IsSBbR/ZKNZDwtSXu5BVpYqJB87/zkpsDXlyM7HGVj/
n5cX8SgBrVcUpRt/ynf46F0s5ufRGcOq6+K7GJoCMpTW/q+Zp9iPzl5BHPwUSVVDQ/Gg8qQ2QCXF
allZbUwBebI71P0ozyKsOYPvs5ASwp9OBVFZwbN3KFAZLMEM8FP2tp/0S+wYkmxsV22uj5zn16f2
bluJFc5RmnRFrtiboPgClqswpmBf5fIIQtlGnoUsmbhUO1ezRCHT6/7iUpH/6VZI0K/EyZf/VRU6
kltNyt3eSFMyx4K7NoFx1DEBOOMW19IgjT1suV+Hb2DyJlUVSi1WQ+T50GKfi/S12E8dKfZ6MJRw
YrsQzsez1/MdGtK2DIGcvo389gNv72I/O0svYCzcTWO8vpYH7VBPWevf5OvQFVT4/0AvcZhwdVEi
wFQEK0e7REMfl7rf5BYc5Q+ZTxkrRmDigQ8TqdfZtWtJeUmh9zuHK8CeLA5kSp8wud686JWj+F1z
b/Q0bVzz2rwFDLdEksvuwh6qILMouWS2oS/TEHtMK43J/FzHkNhQjTPl1yzgGkA1RdY4kQa0rkYu
LYst7njyPAOzOLil14gyTcIMPuJ1CUu0rrRtxNBXlBAG629lpdY9K5okeus0HTBgtnfk08SwSUeQ
RlRFGsmfOFuUfXZOvGxUjIxelsB8NfttV3l1U0HozoaZzNxZ62+Y8DAdasilSXsil7Q9xZOH/bPC
E7gXLn2sO5XFcHnlMMt8qoVdRc+iErWEK91AhnbN+qk3buDfTWuQ0IijbOkgmMAG9UmhomMISJry
oHEmq78SfAfa4mfO6o0XB8RA2MJEBUzvMJ38+01hGwjfEwKZOccRQmLG+/BYMW19A3RDKN3sID1c
yyP0bKuxjGkVzJIgeKl+XL/gtlYWbugMeybuAabqMh/hIrF/REp12qoZnb/CRGaB045Lr8ii8Fo/
A4PHSLDhTQPfKyErNcXWB1jWGZEgAyWrL9MFBQONgHdqONwD1UJQobBme704LuOXayi/2kQg/8S0
shEWuyqDe1pmHsFXNkBRJymS32xS2VW+Hg0HeYFQYdgkAHjT/qYQC4j0ewUWjpj10cLNe5aPDnbp
/TsCy0P6f1ftek7NSYWDOAVHhUm5xRdlXOxh+bvSupW3rysdrUShvz31+iuZ2EvYEDASAXjjA7XT
3CDeS1YiXG2EB5fSGknPb9PPUhDcQyD7a4csWIPdvPWT2VHqaJI+YLxQ7KDOqFpW3RW3nUvlQbJp
wOYC1qPNdXSEMFVf3gGm+OcPRf04HvEai0cRdXwnGGfEWAjUt8P9Ynjpl3/82lY4myTo/9539kkf
hjM6lHLrMXI1D+IuyeKtyCr7OMf31fBZnrfJTn105Nbgl5er8AER3uXDAdgPi2KWXMICw5tj6P2E
HMQgxdsrVc1WePF/Xdz4MKSDMqgEulsaFdoTadk30qEGaSG4/e2zbqczHwuN493rOZuBk68+aBJi
ISoRvpSB1fotQf620MmOd4U4XUMdBXO+zD+HtLXaYX1itcOBa5TjOQUTNpRashc9QB28pfvFI4GC
6AWFSxvv0pfXBVe/x48Vn8phWv2j5RrcdPpsOC/EChw5fnmqClFJlh4RqeWn7RaiV+3uxL8yfkP4
LiDQS1AG7Hz91awdwYCzUmZ3HTq+qh1VICEi6mUFpMYwNDBGpZWE2Zy8ZXrghZvHnncqHf1PH9nY
GVm0+/HeF5oliLpnjThfr/cn9eD77n1b8psJVfenCydmw1N/Mu74WhY8gTUSLc4h/t63Y35/MB2/
ey3gtEecQI7XfGRPapNWMRLREr3hZ/SDVWyBqEG0sSpYdywuzroDW9yIO8KNxZJzGHE2U5fGOU09
U9xl08f4eyF9w5UnOKWH36C/NOi2Tv7x7WhhGzrSCSCC6GRpnyY8yAScfWab+jIGpLhYUxmKElxQ
b9qiY+Zl+niFEU+DUQjarBEc28v3v2joLzEGJnxIjY7ZE2+kU8zdP12fSCdqLykwnv1Ru3wpkTh2
cRbltpWD+a3rTsT3CXalpXRcV8fG/2ar0IsrpqG4Z8r00XeLhrBuu0Bk9xtgzBtY2sVJz0hPllyO
HXHeeKogwhodmODGU9jxgDEIQj7JMYQJtEPxubwrMl5yDzONzFH4JspR8phqTGMAIYyak5xJ4sIH
E/fucoxZpi3sJeeUzDupwC41PTbyagvEcaUudU3m14I/6iA93SxiomH3w3EeLRPwaT3hf7+BNbkh
xHLvX8Dyj5BgN55lbOc6UOdueH+1MeYQrs1TkuEGLfW/MVuhQj739zMwLrfQz9mOSQ8aQITbw6VJ
eOi2mCCWZZtKAKUYdySdI80hdfDB3oV4wdMWG6P//9UJcxniEjQQVlEloBTf6EHxCi9+kxvA7TEg
edm+svfoQ4S0R3oLR/R3NXlKhvqrnMBvg+xjaNtrB/UG1oBKqIZolsEbySyFU9Bj6+vExspsR0TO
5a1sUl/rK62o8SckJ4GNGy2rWypV8rzDJGkgycRke6xBpyYpBBHSTMRuksfAiz79hhm31LGt4DyD
SAZ0oVfUx9pcmVp3Yl9pFrBNV74lgPS7voHC1H/mVEeJsMY5s/QaJE5htWnIjKdVZiHmWBuLBDRp
bhHpmmDAahCNsnNHzZpQKiKapPOswmjLa5bifM7etrHuwF1UIR18NIjikrH0YL4mnR2yVErWPh/g
3aRvA1H75RpAI6uT/ljVh8lcCj8eVktLXspY2TxkKlPjMJap+Xfx9Kd+FdfNbRDNfNhqB4zqA58F
NSRSTwst5vJlx17NUCoG5mYCgEnQM+ZCVqHW/84FRrTB7H6eZnsKd9E8Ent0495ETt7+hG6uGnt5
3ExdzKC32HxXafTwoslbgdI7RDuvjOceR3el8hxbJBcigX4SJV/l2mEmmHan/JAIBNmrGWx5pNfy
PY6uXaLne8l2T7MwookaeiV3dS5N6dzV6Th1vhU8Nvb50vlUlUnN31ZmJitDurgjvZLYqmH/qWqj
9qE95jxF+JJ4zFZVFz6QptjT45mAwp+g3IoAPTx5gpoW189Yr71msWA/j2ESVxpAC/FBJfzubP8I
isf3MDoVwEiHuIAngkno3B1Td+NjsgWq42GblA18a2j/W/ZJxHZi6j5PWzvrg+NDtudY9rRby25k
jpZvx74DHPotywfSAaPkNOC5INVw0fwmSaL6EhyQi9hLqPg/G91il0fREB1MPmjEBpavKo+jGckL
xzjgCuQWgJgx9HXUm2M6wxK4lQQVqa0hyBDT7tCHJxi85jFXUC+K9ua5bhqsY61P/tlkSfNCZFDo
a38lWBKQO6JFFGTqjoxS9H5SLLxqNJmZ2tex7p5kxre6HJLHEbeoW4UnXPduT1sn955Qtak3vRRm
kGuo4AYPnYbpskYNuH82LQ5FotiARwjL36Dr4r2oz26dLRDTcIN02lYCzYCsbXGuCsZjDaaR+sXl
XNen2nh7xbfsucOWfmVLdpXpcCr/r7IpMImDiFJwhUuk0FLqvxxqoTjg1X6lPNxZaXfGaZlgNeei
wX06vPgy3i6PPweapnyopucDBnVe217jDsNRZVRPg6L2Rw3xAMhr0Rbd4loFtMNTTsUPR8qlko8n
tawymdJjXt9FHGxwNF0FPMdJ5ryQKynfWnIsuFwf/JE4iYWI3LsQGy9Nre2g1XLXHpjff3WCYIjx
LBCdkATPoD+oQ8aclQip3jmp1rCcZ59iSsLPzhdfHYBmS8livLN+1rNRgW6NrN3Pe78maMIGV+jH
yVm0oLbCA/r6TtyfCl73TdZly9N5vB1mAjZDF5yKNor6kPdMZmlMxJaeJLSQYOw+6NIQ06vy3mKy
9hvSlWOo3l+/LYlS1wZrBrx3+VQ2cHs2WL4YnlQVUfbi1wJFZl5YfnVhbLv/7tDUOAcA7PjDjRVu
oQOTq9yy5JDK2xzw0fKy6Fsqg4lv9QtSIXBggXVXFP/KEMVaJHxXjJGpqE7afzjMkSDcC83KysWs
TqvKmwcDUDjbTD9DA1cXxKOTXO7/AfH5+nncrjXpzjiTAhAjIOAANmUYfjMJ0IWTr0Dq3COKYCVt
DkGsjBJZkkL0r/nvBzvFChXI+8TvSGV1lOyzqZe/q+ZFeDFhvaZ9jKLmjRBxHgv+tfD+iOJfqA0P
nlGccic8sGKifo8zgon2J0nvAKIVUcIza08Ap/FtfAb2j2lHJh78VmqUex/F4u7+TLOpLlj+30eA
L3GtSGmCfYHsq6hvfDOTZxIswXcK0+oGPnJN4J/kWzuqDXd6KvZtlNzSOBcvbwjfOWlgBgCm/itp
a6PLI2yby+/2O7tUt+4QKKfxr0hHnFtQbB/UsgGiBIaglPE1kPoNb3n6ayJokx779/nODtfky7yR
d790a827Dh4ZkvlU44DOP2Igd6BEb/xlX4wcAAFRd+5JpkarjPe9VbXShEkaix8WSBhV+L0DwJkK
OAXScP1XoHqGdti6bUaPYIUp3g1OOwUOv36lpzfB9YAGfw7FtRgUQ1pdgrjo0jQN0KaCclUcHThi
zy+Uzw9dA7GE3aA36X7MDFgAUqQE5ApKF+971wIe5u1pzDQ21sHMtJlzaqgm7GntZrV44PwZxEv2
Rp0uV6DSoEnKp0me5d9MDalBNp4DthnW7xJ9252ZiCy3beF3uumrWAlItBHgbWHla8Xj2sVTraSh
j8SfaTe3c+BLJXdIaU9pTeNjlxa9X6f98N9mEuFwEzzHNW2LcbpZhmFoi8SHifCs8zH5ASq9DMLn
9YBn1t+JX6/UOv3sRADjKRbJooNXoZUQ1iwNc4OkGp22kX7A8jRIlB/tldf/LVqv8B97jcjfDGxi
O5QYOicqg6okpa0WVO9Taf1rnBnjnlLEOVlxEeMKn5cyAh1WNJJy10BhK6TlWN8xbxYm134Vv153
2SNqQgZllaBCKXvC7CjVHhJ/XNrC/1weQfAFucQL5a10cZjKk7kP5zBJnHLsdIBLKKS9Pjm3zcv8
4h6nXs3x4Pl+T37CFV1sw58WUSh5j95QhtsbM80S+kqLP7kB5zBvilLtAo1owbtAQ5JB77JB07vn
MKjBl4HSaVlmRE9l4LeEiV1tou9i0eNxngRt/fWbfBSuhZRrq2aXNmU1SLRedRuWrjKTkujyRVa7
l0ofgSChNB7RdjASNqRIya1Xj8g+86KnJLOUzRL2oRWJDjQTm5gkRRKKo1DgoKykMwgjb/8fLfhM
LjrtZBHmGikdwxd8pD8VUH+KhMHGAmOdfr0NVgURfyHruFAQzVLM+Jra6FylrdAVu40cliMd7yZd
T6rzFlcYzsCEt77ODTTfbZph5MUCSRXLNDY7sNJX/FXvaGbHihJk2VhAKYS2+btvFrmnM3jT+3xg
7VWDRgAt/8IcZJQMMRlc7aMzutDZxcZDqN4NEH7lb05Z4+L2/iPgUTV25zucEnnkVoEGWtbdSAlB
IE82HJ16t8oadAkYJN2iE6ayt+QxBn0gDbQLbhBPVTX7agQzBey7fnjoWlvnOIKYicIeyp2V1gMM
LUMoh9eEPdZaTzyC/vToswKYss7JCy7q5tdxpzFZPz4RXcxP22u+pOwkW435rE9HdLshckhswDwr
fbZ0j9fiZJU0Npvyv22vF1UjFvc6G4NzDZiJo/4zRRFKSxDhSHk/M0BwgJe68U6nWHAiexS8E7YL
I2zhKzhSpJg4PkYNWlEOowkre61fOLZpVyaS2MHO6PvS7nHiiRC26uW2AgA2WZQo0ph4r6xrtEu6
FnfC9xDEBY+cyRx48BEE8O1JstKaEDhVP/lkU2NC89ivGhCMxiXI6wqmrxcrKDVCiTKVhHGm/kkT
NSABqctDXnKpR0c05BOywhjEie1GU85MLgFM7SpNvbz4NToSEigFp7D/1fv4ZHvJBdiHehqdI2xY
lCxi/70TxF5+qXCNQ7BOMcALUtPRYd/9ID1rNyWTAKvBnwUOnZGyGehgFNbFkZBH0Zc5pag5BpAr
Ki1OExoQQXsqnF62UEAMl4xUlA9FHB27j+NAHzNJAZvSjqQ26OS60AOIAuCY4ns+SvMqrRjPIbrf
oPuIwiU/iiRUluz0FEIhtGjA5bQ3VoPHhBXQUXsCKGvH8jPrJXnSPQ4YjzbfYt+EhKqsiDnoC32C
uGDWc6EWL7a4rnqiQF4I26oDNAMtLA+57dyNPQn62oj6Firwaj98/zm0RAlE5npeECVVtNzG1FD7
O0FcEyICKOepw1s+3F3xeCrbY3Iis9J9mR6A5ETWNWSqkgUwYKSAzopbLMZCqhqOGY1udNZ4hR2b
5Ecn0icGTzCm/3czQCvdhfffcMGTwxWeZwurXFGZPpuMbfBJ2KFfXue1Q3oeKR1OxQyIFkbECWs8
oyH/HEASWPAKVgfnEGd+AangWB2/ld1RsdKyQ7nI+B5v7MZv9Xb7L3l1Clv7SqhCjsWaichwLUE2
WURGYSDOTWl1ptv2SybuWYeHOSwuVvv4D5TfXun0bDvKtpLF0CdPWWy6zPuy6LXUvG/s6LZktt2u
MnntiZ0DEX8WGP8eemh4fR3PxrrbHsuuMNIf/Hs7vZlJTfBg61aC2yU3DGHNxGwSwSnVSNsLQX0t
dWt1Q8zEuF/w8TomSVO5ICFYwMd4qEp5iid3hC0lTRGnJ7tOAq629v/h1liCc1+V3e3bKsuv3+y1
M0XxszdPGt/S5swKs7oNhrLVeP+ObZHToqXt2pdLKE1GsQy9jiEuoTc3c2mLoFaAOfDTRciPVx1E
GQcdvM9RuMfstIwbS41ueC6N7MLsO+CxbCyISOmxJ1SjcFBLemDwPFQc8bFS3NeazpvNFaZ4B8+g
+EXXbvv3oraxBDpN1wubicb2LTQE95iA6iyAuoMhnpJpUHK/PL/QhXN7ZsGXs6Sjtnf/L1SL7Km5
RMmdLCUScdmh0d48n61g7lhZvtCbi689wrPHW0BEZl7OAdZzkaJQaMgc9muHzLvLmYT1oeCyImuh
crNAdSroo23UF8m69Q7NpOX+U15S+EId2wtfncfU/n/AITqXMUDOrXO1Z1kpk9tBJpqGi9Cu1xYl
8WAXYdI2aP3y4MToNB50zSYG/zsQ/aThSlw/0SqwD2M6UfokXlOLjKs7eYAyJ+7jDisTATRl+VWw
TNFTp/SSoaVKJ/jjB5cryIl8GBroE/ITJAKy0vYGS4HBKrhn5nop3lGIVE18iHQcc2SYp7U5X/xe
iSpRXF8xpR/PyVddUghkKNWjcy/fiivDnRc16z70KEgT7axFgHhA8+MemYgz3WRfYdTBxlG7VCVH
5uDYde2hMGptiFlc8BDkJnLgcQwuFBNVSI38UsSJw4HEpAun1uUTid4yS0lUt5kDsbXXLUoF2TeJ
SEkSnQmhMm1KJPZ6yOyRl2EXrTZQYouLbXIwRwqPcUSSG8UPj37atuOAJRsXuGA/+J32pOgtbkUR
ScTt6GsZPwDkzxpl57pk13jVwr8Y88HwwIYHGjU3jPBy7fih6Xc9KRa97ja3EzdupP2gRLq+IHJJ
GAXbhL1oVY/MXyBo8hWHLLuHl/CnrjkZhZGkd69EwLs8lwIWoPSi9YEFDwjBNO1/ZzMYsRBgiiGe
duHoBaItH+1zsG4j+ViLSUSdxyBQ1E32ul9y8cLakBX1Ujs7Kg/CWqDernyW71HsM/PwYKsDv9Qp
L9mwPkc1/X7blmUU/aei0aygleDlIZ5oXTvqb9IaxqAVBDBV3FpwRhf60UJsDZ2k9YdUGwMfxpMz
TnljI4l969J8Ql7nbeOJyNXQYUWCNMNgeTIINa4ng+FfqAN0NSdHzQbg0vQDNRA4ormlN/zAoAto
/STjrwdYo8jHNs9Qz43Wv0CNXOfhr3/8nvNbCXZANrGwMu9uUxGbilMur4AdVxZlCnWtXhjehJdG
6EH0KQYN7i8g7yj4rFYaYP9AIgBCsF5OBnrBfU9DfS3XcPuHfq5pIfuPdKQmdF/AN6ZgkPw2ZA0i
lvST4mHzbyb8Mh6rFhCVP9wcZd+g0RAueZAbTxDYlRJmhkWRFAXd2bW3yarSzb4iu/o45qtA65s4
SAVtLOH6gZKafMVgq0i5oXHsEbvw85WgIdmMLDFz6i2sfP7Dmq+PWnEKgnXViF4fFAeNMAO2gLr1
SIhaeOVxmQY1LcWdeS5W8dwb9emytRwMtnPkt75Lbw2/bOxTAOuwGRaGVCdweIspUXsZ5eYujsec
tdSAtJ0AqUuqiD9z2womkPRp6jo97rojbnHwZRSVeu3Z98nuqmLUA0Xd91stk5yV/8cnshTLvc5z
E+V700d/dsk7FNRfZ39sh3z/47Rd8LLklUpa3RBqd2CISMyIIbOw/nRu+CQU0fgEEIpkD2Ce64T1
gaAryhmDXWBGZl9v8MH05ZJSFmv/MBLydZv5KP15OvyEHoxPyIW9qaci8EAs41nSnCSwdKmnSX8X
UMlghEo+3ky1cruSjRuyinhp6e5CLrSs8OW5b7f7XG2YWcYktQARuNIAqc7yNDvVD/mdh8EbnqiW
DfuYPh9JCqdvpOWIDbAbrQF9i7RMXSGJh6RTLEwNBsz7sx2Fyg7U1m1Gx09reX7GcvNMMRZYPI7S
Ad22gdrVysb8x9U6Ao3c586TxoM7Ebu9ZcOBfZ1nuGNdM7yGM/8foDJoUysilXL+EVPJ3oNO6Hqf
tYBQdFbvkpnizQGppR43mQiWGjvMOCNH6Xp6VWduk9fXf818gx4aX9MLQyD88TXCNEuoQJThbb1Z
TKTzGCeFULp7Gr8BGZvCNyBS10m03syIOI+2JKETVhswIfbbHW9KXJNxII60/cr+Innlnw4BoxXT
OQ8spql0EJRYYBMA07rnSxAfW6pAveP0CQlkyix1bdyZafOVc2EkbE/Dcyg7zr2FswDn+lwjk5nH
7pVfohcntHYYYw5CtvjsJQt+LI3mlutQ9L5viB39JP4dSropwDhtnQoixrIxKxtCfF0787JCQJxR
9q8z5IEEikyNBeIXvhLUmq1KB3YlUBsjjoSKZaG2OIKJfoZ7poF0sgGoRmJFiZv7/s3u4pcSV7dD
e4azEYWsJ/CNc49aMPNW4EFXblgMyhqr4/xeW4RkJYUqqw1ei0zst3gnbL619/9Mq/znPCPS7lc1
OrI64BkWsqrGUdTQIvuTXwTxRbvHvlonRj7BlYI2LxlBd617DP1zf4OntuOAn+UKsBUyLwyzPL+E
aG1canPWPCXj0mKYq3xxw41pKczDs8XEL2KrZ+ii0riSN9W0OXrMWtjlAgK21uJdqPZyQLzZ0Evj
vkfjaBpvSJc+3p1r5TW15GN6OEq9acDU33h2DV6QfactYtiyHdfD7wZbV+JVVINzfuvBFUWDf55h
PK6WpA9UK+pUhl10ZErnnpn+zmmVZuQH9qtmG0o9P8CM8gYOuv5cDbiwbv7EiipoWwawvrECa2mA
V/eNlmruVG8ekjFzPHsK+6AA9y79zHxvGHB1twDwJ8TeDyHkt3/U0kCQwJdvj5YbeMzKEMl9o6lQ
skQQVE1dphqqyJQumX3L31odb2ZSaZlMkWCeuv0vzhUq9QsIicOyL4dOVgAxvU5rHP3xv4RYDnVJ
QBEb/lQMriLZjJ0r/mJPhp9T18LQ3j/C1mnVzz30X4ilHws7HZ0a3cThRVvygFSFM6hR3eDvD2m5
UY9Z0VtqkX3CHjKKsM4+K7f9FBf14lwJ7wZLA+aTvtHvgrn0d8GG+lz/Hq0OurdvVtyV8asFSOTI
PH3EoeER8vF/eQBLx72rCyEgm1c/9dDtkdqIZRCwEeAZoWVXmbkTIvFFQCNkDPvpqgFj7Fqw/jBg
GFItZmLjdAj1byx0EaKPFoVCZ+kAVowPkPqIWFjES4tCw26+Iw9epUj/60FWQ7w57mDhyb1V131I
2WAdu6Nn/Xgk6k8hNS7hf6KAzvBJsKsCqh0QuGUJP/d/c5Y53H3AqIIxSV5bYDaSCCP6YclpgEGv
7aION7GXIMpHjj9lVQCKIZlA8h4jr34UV8hso1xLHVBnQ2nUpccYgTPi19y3k3296mZK/69vWmFF
jNtCZbDKu+mP53+eiDYkBNMnt7gqa1yvEAikx2kvw8U7YngmML2jak+6zTbuVo7OVNmPkzYkQO7g
AR3pbV5Px5nlYhzniu3HU/d80zWClUYfDzLT6wvtv5xCYksRenIaYzGT9L8pJguZ3QsZJAyhUqtm
19zoJUTw13025iwgHFMA8bXmkdpKCM0d9YzmX1JjOxIvGFWvBkFVg83acuNnjEvlf2J+jPVOs319
mX+BncuXXiKQzmgv9csE6zOggk1oCAF32+UaH1lmCVvy9ogMA+GgNm5oJW30rDV5xWkDcjufxQZL
O+yYnCgLHr4ZyxHbGSE1oXtlLuLrhCbe3KNA3T4Pzs2wgN6xQBvjgPv6hN4Dq8WMa1Y7yLWQIr7R
YF5p7htDPGgHM646QX7R1J7SQWeE4M2PbtTR92GCMxyJ0nJvxGdZMFgl0lgHv10o++LROzbBonc+
oAK0m5i320CiNZKvds5RSblVHJ8LaM8alfWCuE78advMZ2SoThNGDYlI5nUE2Nw22NVVExJ1HTxj
pQmayASkhivMdWc4MmuXdvHnZ9Ph3Z/pJ7jpWmDQGxCqpIGi2D3w6XeWkpp7gU49O9JIfaCnQHX6
AoW5n5JCe9WhcVbO/YsbByZJjlx458ayP+cHHLDvgrk08xncq1HMgbck8vB2F8TZMCzKVI9FazIn
Hx22Jl1NzPlcfwUWGV5H8tBdSx7jD+D5WXVNIC253lBlhUX9wGNmofiFfog1bYhIATBPB1c8zXko
wfCSBlqGfA2AHkicdEkuqpT4+wY2+OGQTj5+9ec4h9Fj9CkpI0G6YfpAES1FGJDUt5OEpO64xRpv
oIyNRldCiTEF0zyjYaqpmYoyzbSBHE875sU1WibZI7V/IqQjmaY1OIxG/XwCBb1jhhRd3KPURUUn
5yZ7bcQmAoXyUnGt8DJz1HVDS5GoiCEBFKKVuH6JC/SUdc+abpaJhqAsaYP8gyns21HRadSHgURs
zdQoXvorXknl7I2xfMcuEciMeRXkmGCy17iizkYUcAYL2wvfbxin66macwQsk093prnnEd32WbYb
HLPwJsre1QlbcY/N5Xt2JvbA8znhDfP7DHA181jFq2Q7BiMi1GozdYe6l6DWzVwYJhlqvpaLh/XI
waRHONpFpgMXQOf2uJWyFGpIk+hUaT+9IWkXppJtKV/MyPxT+uIzIOy3m7suMMXWkHViZyXohilh
aNmftubzSnyQPds107XEslw7wMz5uSV2CaaR3pft532ptcIiRAZqOAN+FiuKqRmsLyzhLkAhnp27
dyRZ9GrV0RKUUmwU/96YUdiSfuOu+KD/FwbBrYMdt5CqZcLBobgldFzpiHwBjZtubQfzWBfuoEX2
dW4DGBcKabgx9wp7d+JmyRapwDmNiUgaFmIlWnuxJFRf5E9QjDLkrvovXpibAtwyGmEjCt5uAWwj
g075BgEA9qHebS7ysToM8zivzBeA0dkxDaBdcYFsk7qWd6Dfp5N8RqD/OCzARhTuC+0F51fUWBXA
bNciW8SMwmZXVIcOhWHEkj9E0ZVCLEQ2vaUC7EQ2XgN/H0UEGf/3BjDSC+oYvQqBiS0LRF3xHHzo
USnCybWxB2/HAL+Xl3vAbxkJ7awx3u8Uqlb2Nq3AWsuFr9KPM/2k1b7ghuVqQQ1Qjoi0GcCej/Ck
XfEV/XN3FZcwB2/XbllTx9H4Xx7jMN1cMvv+8SG9ZlLpjXKUjUkNtr4hrLkRZmrrDU5IHtI1bIVC
c/QZT0fwPbF9F+5EuCyyzAJEMq2xN8CRRrhSozoVlQ7hoWnXA2T0sRuiCBx49KCcTjv7fRU3XvDs
/CGSNeZ5Z4QcdVVN367FqVaJauhWOb9vHjTr5D5s84gq4WzeQiXPlVstIKil3f2MnFW8JGAs95Q2
HRswCrQs7zUUX7BAN8x4Z8US36XO739N4EesIlcxNjEFR1Npnexb4zwZIASwKoaubjhlrOlJ35Z1
LLPGu8ZZHBJe/xHryToS6DatLdeT25AyfDy30mo44DSvEV7tldm8L0B+ZZ9EThbsqjQPsdlkMntc
sVUNY731zd5EfbcpQEwLwgnvkgpgLLHFNeBZi+HMiOah1U3BqJyyGq9XFxZKxC9f1k4SeS9qnzQm
h1WGi7HlPLhHZLCVLJKvbMPef00g3/FU/73XHCCXQ1xOlnCNEYxr6MNcnIegbL+pSqwLAiI4i/lo
TfZ3QUvIZODX0nkuUOQ2WYYCCB27mVcmDg5eoGazcTO+WlynQsXszZMVpAIgRSf5AxcPUsIGjn+O
oBmmAi3XUsDvRRuVuNEfbfcnWDsdmB7ImNRA8v0JAeWqMtUP5E354/q3vJa1NIaMXUT93AepJCIS
S72ZX8ViOs05W4QvR2/63kzjCiYmig7nB2YC+zW6TvQJY+LRAhj1z8mo3UwF5KkVnNnIpFdWUobA
9NPmr8VGmK96SBYUBK4a725Vxrajen7HOo7MdJQ5sRLI7jvhEbEhxOmvV5WhVttp5m7WLrbJCm3r
2P9hegUDPn159NZSMv0+eOyY7+gRtrTvYMHXotCH5HS/ivzywZK3y2jbf7QjqCVHlgjaKcv3kzq2
uT5Rp1wwJlwPyAGHzNdJ+9qAvuDP1xK8W50Eprq4FdLsvV+Tq1xMkEtIgzjDzuohg32LQ+74mbG4
tMnyODVqBp21nG7z/cFkALgVzbZE2xRFWCJCDOs1GjgArTCRbYDkE3wALKD7/tW76xBosWHyZAhB
MULnWjdPD+/sG6iTp8IORBAucql/muU7N9GuEiXGkc7VCKY6n9TMLoJlBy5wNstUfE+MHNFJ29h7
N7WqpbrrmcZOoEaQasd9Bvmqv3Fnd3o8aAW1jcTViVBm1+PYUcv02Zr9z/iBqZXFNmivDbneHtbs
4xbPu6lhIDQckyMtla7QWd4yW5vKgSRNQXGCxgFszGBK3cN0t7KUYQxZnSBw14Y6Id8U3D4YtcuX
Yj9WAywQtPMzv4bKcC2OSKQK1D6+ShtR0hURG6XRdzTBBmHWatxHZOQ2RLysaVdY/AUeIEkbhrCA
E49QPBXnW9ULEYzJXlD07Z2SBtRNLZCEsaZ6fjP+8gjteOLOkh47HiHM8xeraMvOR8E4LsXe45wF
8Nz2OQUcAcsfoHvGQ8WwDYqA8yiZJ/AwZkw8Z/bwbyVliF+O3GFK4z8D0e3Wtn68DlHuk5xMEVJj
j8Z4+s2LqQNs7Ll3Mi+OWGpC1gHdH2GmBGWIDwVLq1MoPYixVRUwARBNOD31ToQpZ5fEFTJ93wwc
7oNyKns65zz4TzJH80ocpx+yGQo3/5827SvAivOatBMQ9H/ilYqd9DhGHULHYHk7ku8rRNItEwBA
vnnfD0ljVP/NRtennPsXImvbRzmyDgifn8EZFdIuTIofb0MfwbY0gYz6/tSmWUtA+556FvV9oNSC
z4f/j3r0B0cX3srmwlcRrKP1GqFN/GjVKGyCdeXjtV27wKDZEL998+c/n+WhKH3A9hQjMM37PJrF
ITt8u+XhEUTfAHP6fUJjtDHudmA/ywd/la9bDDWeJTUzW3kycGdJ0rDbMCVCN/fZC21fcN7SSotF
xE0zWqUEsf19rwDhmdCmWhdPI5CHHvKd/m994zlBJ3E2xwYZCeGjJCQo8u2ns9BOGBVtk15KaKQ0
qJvsWB88gcmheeTOCMDF0v3+C/yO0MLXAi3d23vCRS/fQPQ2fqXwy2wYdLKUfHD1HpxmsfTEepCL
h8vZZLr4buClxSEDmg2L2i0H7yaCidtrzO60444HqNxY36bPsOuPB8CGghwberpAV+YqPmxT5Kts
1ouei8+8LhjGlG7Oy0cTxKgR8MNuAls4J/XiIsUOnRUHYL7uRiAtFsib53xaJQVUpsergpYCg3O8
hA4R19AXR+p/2jiK3ImFf9OYDqr0K9IklgpxM0uEG4viWssTIu+usCcGoHD1GBuPc2/0YbunnVan
68BY6GRX9Ak3nKK+iYHOR/OOGivXaipQke/ZWe9Ba4rKjDSjHUvqRpwHCuVSY+abNYK6Bpeg6owL
1SIutO3lxd0JqeYtxEIFyBMbPdNG4BdYyuO73mjlzPtjN5euMYrg8c1ZuW4lkGuFyKVXnWnMkU1s
oGiRxAOhxg4Iasa4lQIxSd5G5R7QHU9/NMQRDLcfEDzMw4hzK3T2GCFYTQaskNAuHlIALLXYua44
dXswuVi61Sb7H1KHLu4P/7y7ouNlVHLJQRM0YD9xFDRmoNgaUvRAnC8ywsFu+1Q6Rzjxa1aEnHDS
a2yWOUSSx8SDuAjp+Qm1f9M8/pC6LbD6hAqxrYyR3yHU9cryCRVgam7CJhkywQ6CE+hXTuS+tVGO
s5iE8iEXv2r3aqbZOgpnw/pPz5nOUU1ewIVMi9KqItgG7Qv9D73QmHz2n0yZUQEE1cZWC7WyNf58
JArvElhMMN8V+WoZlLZCAv5BWB0mPSEBMA8LDKjTJJeIj/4I+6acXOi3D3cBF7QB5gIyvld0Iy0f
JZUTV8DjdQQ19QOUy6a2YfQEkB90wg/BBczWaTJyhAzkyrP2YUxo1ZlXQIRE6TgRdwqorf6hLp6z
S4NHrPABkWIixJf/DRmDv9BzlpWuNAssDqHbjKCmDHyT/CNIaAE5JcB9EaJwr+FXQJ7LtkSx5stc
MYRzgXEW7SIkfrY68gMNyqoRdtTu7mWZTbd/gktI3ZEbKd2cyfDkO2pBtOXw/1VnsrRcfirhit9g
rBpiubim2ckmcjaNVumSRS4g50rrGPPV6LYV6Nn+thJkKfW8ELRyq5QGJ2bgt2J0E3Ha8TbZpkRO
TlZ0D/pp6pcz72oyJmXtuKJbrvbtDzfdG81mnyvRV93/HxaSm4E4im6rLs1vc3YMIQUJDOGRVs8m
sCoRxeZXg2mZan5UZub8xcXGjMcdKJkPLMeS8wZBkjKEube/OmHDa/uopuO3Z8YqQYl4+MVLET/l
1/TTE3U3o4JI1woZ2xaTklWspTeSPn8otatcXwgkyJZlE1+jeMQAbib8CYa1ntGOsexKI+W3jzCc
+lvvZ14JW3DTeN/Mv895DsA+kWA+rifPRQS5N0d9rLAa/Sd2yZhhlz3LepzlX/qh+lEy5uD+sjKP
XVPRevQfDbL/1shGXnrV7pCMR8+EtL9+BZTK/TE3jO9uci+qIBcocckOsEDOKaC3w9oBluSeWsX+
O4gMc7O7RdJ4dlwLOmmMV3yNPXe06o+mXbKdhsI82ISOFHYF8THtmZmnLadVXogNchPzSiCIatKL
tVf9Q9rEYQpxF3MqIJlbyru4UXa+sNbv1ez0U6uMMuaPZnn8+RS6hUbcatwMoqUk2LiZ+TzWXv4/
tEHj14SQhQmC50DgeBtZZ0vzECGykcpI02U1mGxRTvwFBEnt9LIgaRXqMG97mjPvdWUDDMDL4RYo
w34JQDo2fSMTEPfuMH437RcrSiBFKQ2V05cpFhKsQbG6b+HN1X0pKQozWKPCUoq2ikwV6T2xrqhm
gOKVc4EvufbGOKqmjBhVfNpY7H0YB5f1rUJn2UwUPo7EJA27FXUuJVIbe3dJwRz8D3/qhgjU9nZO
ziyzTYjiO8SoOtlJ2vVXyxsSsTa4pdLaFFm5um9oWhgQodXkXKsWnv14su1H1VB/d9OV6e5/8Q4E
b2u0qmA/KACcGodP83Yb881Yt8Q6cD6RfhuYHT7JxjOtDtdwNRLU5YYfRjskxYybJBbL41yMEZAv
56nvH16sxILyXGAB7stzwLBKol9QiTRUxouNfndacnbUWePMordc8TMkBjavFbXTP98TluaAQ9Gk
aeO8JR0is68l5Qit85rLOtFxdr7J6ZMbcPifzoK1yjWoY0cP2HTGgrxxsL0d4Dk+I1WfTI1P8L9g
NBFabL06gJuuL/tSLs4/ikf+/rjsWfePEYy792kH7XqRIfFmTUsOcfqHF0VaPdDQFtxO+J2R3EL+
ki7zXIGEYbLm6Nc1Ev5ZpwWCq8iVrtxqJlQxJ7dawC5iXCoWz4xJB5SHh1pA+LGvbhwotr4HNkzQ
0idhflT/UZT9uf04Pu9tDF+RGo/zNnUdqvNw9U70USyN2MA5lZh4x/WLN//XQECv1hKbNwNdb1jl
fh5zmqiZJ7UvJUq56+5vuA5Iy7YX2iza2oUnIqviUpmCHinbLs7tl1daHzYMxoSMq46+t7C4v0qj
S57Gne7NLP3J6CE7Et/DMXJi8tRGJrW6y/o7KeKJkE0odBxAF/sRBMerDXFXSk8JiShaTOfRyYVn
OBa5beQygXyo5GAxRh1d/yapTjdYOoSpPUm7r4jE72+9p1DAFTf+YneGkUlSoXueowxftb+y9tgL
M1W5wINC0VahZOyX/n/MQX5l4y3wvp5zUE8gijo3YauONbKmoKI3zjsOnykeviiuwTxuX6rydzIb
zuIeIl0zv51/eUJj8pwFgVBmhYYfl0qAAEeSOInFRAUA8dp11J80Y1vSlP0VwJIZn1eJU1rm+sAS
bbLtQjFlsRajPQMzPELdJyDXV2cQAkYXJkWHdfamV5/skk41P+FeQgv8MNU2gUCtzSOR1S3ULMxJ
HnKYNvFQl8jxZ7cXEf3TRjxOPr57KekJc6Ox9JhtIIkxt1Vy1k6U9KstY59C8m8YFl1usDXL03UH
/J+xFdmiBIEcJPfyrZxerJ2Ay+jkkrrXCO1Odfva3oeVgdYR6+VI1pO6BQ77vFtBZsXzaMOWFki9
IL5J7bObt/PphdhiAABTSSpfptblh0RZ6Fvarqu519mnVi3sKiD20PvI0t4Ccjghv0fUFUVqCz4c
bTI7jvDuxHOVzUev1AoSQWAS5zqyVGoSRAHt1r/7QD1YkExW2T0z6wInuzZ6EQksKlairv0heuzE
CUiVM2d/0skRNgIfOrsbWnQGK0Bp3W6f7Cxc9XR1HQErF2W5EzVMIOa+CmHMgaE3W3dwOjXVI3Cb
ubLxp0qn5B9ZABFQJP3Ex72EkHMssaVAm62O/GUxiM1+PMWRMXEG8w0KYcrOSECeJaouBs7VzXsV
lCOGIK7rxmDpGBQS7VRJOwh5CGRXQhzpgtkY8Fyf8rHzig7IXlPizVu8quXtAbcTks1xVuOwrd2X
GLNuMAoF63ID0cO2GKhPQsqhSMDaGZVqIzNbTZ618/qSy2XiI0QMgso3nT7ihgg3izGuobqs/gmc
KdZ7zyOF0bD1lSU7/Rtt2A7TGtYc0LVNrl6ALtywI8aPvaX/uoz3FuS9ZPpTeosiKvUi5qbhbZFg
qSFIK14KWpr0nmO4lPL0QN9taLtv40uSBNXS+JDkohDrosoUNBbijVJeHh3RgsXWoO2bsxcGrJ5g
CiSPfj7sH4AFKnL5VRZo64ovP1sLeo6WxZc3dkGHIzpehH7F0sIpRzeAJvEOFcZzw5i4w7gTmzfw
Kw8EDygj65AosvVEIdN8C/DsCvRBLfmFCkT6S6K+mZYRZsLG2rf3xHFiIID1J3Ikwzmii9zNx/4C
8nnbLCUJUYkyzSjMjF/k1D06bCBfbh+FVWIpfiZr/SUxrR2vZybNEYey9zWAKSQhFuSfWa9pw4o5
lkSf4R7SE7Ah2L2SNNqtGKHdNtVoaBKytuzWfGKXQ2fryO0td3xL9ACPxQdDOb+8rh7MqQCIu5Uh
y4914ddUBgKPG9bbLsrY/JDWT6AozGm0Ah4NI0jXl6hxmpAYmeWwj+DJCOaohlRKTZ5Xg3s9Tbzs
iQDgqp7l2pSihkwYUNP23ZYyZkJBClOhYeW/6NoMqD3rE4Yj1A/gLWvmYFUyKhcVWuSigXhkM9Dv
iA38bsLrvqef2v0rdd+liFuqQZRCE/GeRhzs49uJBiWOJ4b/QwEOFnLgbO2CY4P7misths87wKpw
OSEeLLRJ2Q01eV2II86SakWBs/yeawcuyYsmg8a3rmoFhpk6K913hm2zK2xlrkgZFkWy90yxfEfF
L6ZJhcQTYCCFii6MAt+0/TQI8vffVmviZbEWlwCi5eUigOI/8oikMjkkmtgKYrKUddMgm+q6No84
fWY+ocC8n+q9Q9Sm3EyOZzXKrQsM3wF/OdzeSO9GV9K1P98Psx/DjJBCsw4Kp+kzEmlYY8V0X6xV
6RhC6w92p4PrKsDfU8hg/dbUxazfZgTrFPIReGadiVm56LNhtCtFflxs9T7Z0pQ5cDeFOYHXuMET
2mgt2eaE7pa1Y1zWynWH5QfjIJQLgGoHWjWgRsWkmowsF8UyhfFG7pJyQBX8WcpGTpIi4s5u/bYu
X2o28Qo3CQlEL2FTn34K1G9Uh5d/PqSgAwhP+YXE7MgJsBkLdppmZ9Q9SZru0dNjmBG3n8jWEmwf
Rexk97f+1UzraFiCyzZnp8RFpYA9ICmb61A2PW9/mfByPcyEt4OgOv+Sd+ZfcJVW1pIkTwbCYC7O
2LgHgAONFqIzBbbr1Z329GCa6JlmprV2d2toHiiTAxeL7iol6YTyXD8faZYOG5Kz5YtuqSgKOftd
geAVjDNOm3pr2lEgpbQd3S/IjCh3ohZ/jebmQvmJRD9155JcGOd+a91rDkvj+aX9pFJojw3kgku9
0MsaT8PBKT3HwD3N7Q/SkYH9pfZvbZV7GJqRNOP4up88vnTgv5kH9/g2QeX3aFKKNtoxEPI2G/3M
1apgS2pGHVWdikaCEmkoxM+vhynuv2gEmCrY64nsP7bVvVW942WuRVBOQJcSYBW/pjTGU8vW3XpM
9vzyu/jDFCFKzJ8Y+O7ZfMZk1/86a7uN6LluOkMcueh70wJLQmIas3ekYUf5RHrpoHmdKS3Qh4Hl
Nbu0/sA/cvDVGHriVPI0nk3/N0dIh+ZboVR84q3Ypn78bGkR43rWZXLqI9deTXj2oZD6KJINj76h
3yS21gijyR25he123CzJB6oMP1eS6Dz21GCdt2J/HaNpatRP6alV6EVidFR1LWIONZQkQbJqKFqm
OKA4hU3Rdl6Q50wKi17y3sGvuriNY8j7O0A37dV7ZEFLayNkFRB3/51tV/JNSSUSUPVekq1vEx4p
G/0o4rTCO9rPcHT0R5cMylTEOZTxbUcwn8hEl2uF6sIgkbNVDcLscjMEspYx4NfPmRX0Rkq30EYa
ddAaRaO0Sx6mYC8aI0CiTzy8z8D2d8qAjNhV/mgLfk9vpEM5TBOWE+6bADgpP0V38jqYym5FZzf4
KHRKVD4jHRTg9uHLUBCjOP5foNhfyk3fngv3PuJhqf/rsD2T0AoRWXzNtX6ig6CZjqJDIU0PqYsq
g+59YlbxoDARJLwBP4aBn3jhQvN0imaKlXGrX4IXC8GlLhWW+4Gp6zyQEvZTkbB6PVWgkBmv5Bq/
QGOa50DyxPij2axIQpIWP0MLF9klZPAdbXGqEh+eCIRtqnScTtMVkE2AQtvpwuhwkjwOxNNCdjvh
kNK3PW2vnxTx7iLUFBJ3mV0I4y+EBQ0mPWDycbeBCEhQTpyb+FPw9joIrBybAw2YANSNE0x1K31K
pubdENt4e8u4HB1Avh0KL6jdq1elYPym9fQDFo5SGfU2WXxHY3T7JGshLCJ/MK3HQAxFTzkTw292
MwOlRTdss+ggTivaVrazsCsN0rgar9ilQQSZKnZ1shfITwmEd5eGBXpl9abTodT6Z+Vwfllqyng0
9szLo8tBMO2Kgipv86Ciuh4O7KAAg3dmQxgo1puPIOwCFChYs1P+Mb9ys05TN/fNQTDEs4RMVptf
/5+gGiMUqP5a/3Biygjfv1dmeVkoNVlF5WllDYowimVnPq1nUfuE1OL7MGBa/7wFpYFo0qWKw7Mi
fXppP5giP9y6974itsJX/X/7HXs3DgXzOq3WHvqNhSy8ZjAmiQvdqJxB7lcMTrQv8SK/8/TwIVIF
L6M5GFsea/VGb1CEQB2ASGpNv0iyL3TOwAl8kuOOI4z3cBlwmQb9x+48bHDjBXDkvzOo4nZJL2jY
lNxqL3hJ+8J3YZ/50WyAPLiizqCZdYVVqQ5q6LbUK4QPXDehLcDK1FwKqvAOILSh9LHNPGkpND0k
tnJJq5r8/BjonBuxcq7utB4h1Ho0/5SRvSWQ/1JjDi67xEbQA5Lk02a+qF/v+PueO6wwycw7hwFj
oQs/WKCsZwXYtx9qrhyFvsvjOORcNfj3hTUjA0u2tprwFk3IiDWegS6WtpjsANOJeVMRWvSjrgrr
uBC7ipbG31+8ycRRaLTxNVnmGdqkTQxBfK8UHU38C8vlmnVeM46HaD+Upwa+iRVvz2lMm6fFtJ7Z
gKHy/BI4UxBNYC/k2/JTN1vfD9nV4M/1SqtLv5az4pH0pN+zCiy2NIpMsWF3amPlFODKq8G+IMl9
00iJMEKpkuGURVn/wPrc4IBrdzOR09j1oYI7C/cHZl5qZYDkfmF1eLbVSQSkJ8E03DFMsYApAA0J
Tc7ZazuzEKn2ZNFwkrXiL1sPckt2ohyj99qP35eHGBuE1PrsxdzgdZGw8VZ0mOSpJ9EJ76mx2yJE
LDIbojp/MTGTH9S8a1HEVoaEzVfOBYlAyARNREZ/60aQQpKyzok7MusWxMwYMOsRRZbJVnXkwtic
OVP1F3fYlBH/b4YTlqTlu09lKk/nEMreqD8uIsOL4+ojBp005Xkl/SY0euQErXr/CD7qGiddv8Mh
k9bNmJwpXGrzzbMZjZTARcrFcBylJwc6S9zS9mgyiOYNOGaTEuNHOTY5p00FJ2IXLPpql0tO81sW
paRhjiPac4pTEw/62BkcPk48wBcodzBWIhmFeBE3HunFaOqPBkry9ZyiURlPC3wff03S82pgZ78A
aV2bb20PuyvF0TSIXBheyAebebfA5I3ceQKNYczQaZWGtpKCYAAMCZJk/HE8+9DR2UXXvEQqBu1H
xgLE+WXQEeNHIb4pBEXJVC/punZCFp6zXHVifLVilLfcDdPjeR7HpCacLDCIFxC21JhhExuOejO2
+F9lomC6IVT7t/rzrQYw454+i5bG8318M62jfAZJurg5GzDm+g2wrOaNqHL6eHHgac6tiW6rbQ3V
2h+Gu/QFIqsRHrjwiYkH2OXmEc93RLpp3lolQykRnGU/b6py8xcIGZVQvqNagj0U1C0GgEwiwjjK
wvWH6wGIXHjWDM1ZENHKcD3x4ygkYNkFQKPvFb7qxQubG5I6aQhRlxq4XMLEug50mknUesOKKNfA
jA6DKvljfuJW0ux03/D6xsu5gai/u8Iyxc8MDVrRU2kYvFIwvvjed62BtKHfQnQnNxuiOefy9/NV
84RscEu88KtqO8ZqRGVoPZ8i1b9yhQ+AAVltqauqd29o3wGTNBC4s0lhRTpXW2Cif1WXW03CMxnn
KjlXM0322iqUgAAdQ6wLk0+m2P7Tp7MGi0LjpE9C5BU97r7zb1JC4mAmN3GDphyomBHdA/TcHuhX
4NCEZVuzB+4DdVCvgV4crbQljGXoho+QQw5YBmZSXBMlUkX5sKXSUFSBxX4h6BQlFKctaRYn6yhB
bUUYEfrp2s7L/vGybKc8zBWjH5Dj/eLm2pAgL5ryGN3tGMT5AFE6WprWNU39BPmlJXUWx1FYN5gY
mPEcm4hEEhv34Q6FGNWuABZkVELTaP4C0gBg4yGx5iSmeZ+OhVkUA7V0QrJ7djAm6oZPdIiE+wj/
4Gb8t2EftZ/NBeQ93snNd9xC7VQ/2Bzhj+mgQrfoy8mEhbsbdkGtXLS4cXP/rhufy9wyAzZqPh2x
KgC3+hPEoc9ztDdyNa5qPgLsgjOWT3fG+MdAhBmWYIL2ismEUVDP+IMVUrUut6TrRNKVNzHAlRrr
rLwUfBjw7A/wpof1meGoix1uS/i8RIRwq+eR/51sgHahoLuc7MF6Dhs1jnEMTuqAwKkvQvBXQye2
5Dd/zLn0D381gMN3TQhYFGAj7H2ixSjfp+ZJRAuBmxQtEUinXkKak8X7M2Kw9vB6yLBsvPQKjvE8
Wk6v4q0f+5hoZ6F+LvFa4XjMRumWPAeI2xlLSWOHz09eBUt9/F58KTKv68HgpdHKv7gRiQTuz+Ji
ANU2uRo6UXxRxDyUtINMA9Ds2fIfQ34Na6v456kRVZCEezQW/Tr1mpXawcb/aZeIJXgMyxpbKeAX
wQjWxlyUNP+TVj0YCF0FpspyqMKTEFux6Jk4myj2iASNo+p8E7Lj41DL31B2gEeI4aAe9GA2dL3x
nOAP5wbeFcZK5hsZpsj4mKdpG/5IM4BftIB9glQ9xhYeugd8fS2t+PgSdCqb8tYwJ6zEiTdXj9E4
DO9Fd1TDvh1ug3lr8RLi4IuwBM8ltkVo5Lxg14w78afHtGGQpVTrtdRcB4jonAdGSX/Wi6tZhPeX
HLeE0aWqb6UlSzOe+xkiSqF1Wj04YHN32MdR+iBuMNl8ChBkGWtRreXf1of2yEoyfC+J9u62P35Q
bnkJMBKpcdVpVEhV5CIIUVgXgQpOL6uYp7QAnUYWc1LpWELEU+TNYA4l4A4akQrsA9BxfWLWJawh
Rd0FP6CEOQC5SyoJQSu+BqyA1aOrYnomDb1A0sUvSDjHl2njL3SJrOt/JCMy7dL0zJ8yrX9Gpq+q
h97RV3K/GQtuCOTP+KZaNlIW/eqwpTlObYPIo2Bnp50CnggXjbYIz/4/lTMM/TYwgUto0SFzXuqp
XChyIpppe4VYhr0HXu5AJgdlgorB/SW7qcuRKNncXY0ETPnBEa2iXEZfRbDJlr3X/b8uA9LHkHFS
w5CCUNubD4qG3qH7+0vybWq8oSD5aTxRdWUym4p4hW/Rgi4qbwa6X8JZl77mKVIWcecCWeA9r9ka
wKR8u7vkO/vJsdEIR0Ahgx2G8CH+NmqEhRPJX9eix/j2HXKQIjYZLVn3ritcok3FkEW2F29zQ5lU
LaMzuvJEV81XT3YFVBcnbl08nfKKLBoWZmSN7InPEHpWZoa3CV39DNVrz4624NONTYHodlfT4ppA
WS/ejmGQ12u4LTZ1O5vzeFWT6nurcP50zYut+8Rqktb6tp+G0i4fKc/TKKS+UbEyINl+ilYZuwGb
Q6hNi1pee48VTeMcjtz1drTr8W2DfLbK+6v/OBKP75SAIvsQAbjd9qykXV7oQiRupZdyA2l6Jo/+
RyIjnA/iyyIkOAXr2oADfaHVGZsZnYqhEwTZVZx5TVR1c6jbgavzm1ww3mv8YiiN5Gao0AY797TK
7H4ZcMmMeZwt/cRQ4J1ZRigS8GHoOP42WgyANbYzNPXcqtasIkX7xVfcq9JxwazF6D4LXzn12TrU
tMYaVNNICvsKZBoQyFqkqLIprAE9SoIeI27SSi66FuwHd5VK6o08YmI5BF2iUJy3OEyNAuwBTgb+
mmL8ok2VtD0MqIhVbuUOR/uzVC5I7DL1ViFuGLlOOBJvL6wlrvBCYfYHGKfd66HE6HQCX2S70wum
INy7ccFgMVUscPI++Gu/TX/9ji0RqdSwkG9EL7mGEG8qeNzqJJJ3tdfb2NOw+4mYVbZr5H27SfqP
m8KlU1Pr2nx+//2B0UPbUdQy+6Hp4JdrwXG6iZQRlZvJdy1kitf5HEA+77zWMCDVsv1OhUyH1rqh
q4nMuPrG7yfg2Ph4Dl/Qctdd4rch31XdwLqNoTEoNkG1QSPL8s847kq2V9mwAqyXu2oZmdLQkeZ/
TiL5mGeyn6MbBDRSzfK6NKAwh5IQDW23YBDN+ysmfAiEpx+cWwyBKkkY7FetIKHshq7duJIQUMgW
qVPM4hGCyDV8hmmAHaGkXr6JNwUuisCIHisyK5hjotBuFSxZQ6/tkhA3QsyeUEO20wcnKv2cpPLp
FAQuaomsYuVoQuSwoO7kkHvLST5YkbzWKSCdPe4jpiQgsqCQd1zgvcOkYiMvGTqssM5+qotupjHX
1mufsU4zqG+Hlm/ZOjJ8aerJ2lXKG4zeSpZ3w6p9bKuCjQMQBK7/7zxCY+utXzdI4eKZYWh9jAwM
1Bal2bAPj3AdwJoVpFBJU62zAjS+t7kLvMpMI99/JBdebJvguLFeFJnFl8c5+DnFhRAogtee7luh
fQP5EbT+vNhgm1VPEDrUtbXuB1CZo1M4ApkwwCR6k4oy4Zn+reAGoUl3hQUKAiVcmUY17XoD+WKO
+AYRq3NJHh/lWZOv0uu1nK+3Wmh80KC8QdNduLfhpVFWJZ4+z59lLvI4KTl/mu1PkQH/CVB5d5r1
cAVW9jKzJR+lMf8JDqXwLiZh0IacHDyp5Z9jtuLrnsC5XsZQR9J7nkTTkGE3wk9cSMvswrIq1GTw
fuPJqFljm/fhMj6HhUZJSkQy3gCmR6lOm1s/RK6Ja7KADlGr19tIY2177ZCOnWJeCxlNGQSfa17a
hbVAwATirEM7iCHZGB4es6KpeIMinuRvUW4UV00ujYx64iETr5J8rxHUWegDRYQjwAIp7EFK60nn
EsWynmo+RZdjlz5d586TbCFK6xwnh1wlNLs1nZErEBLM4DHEjMDQXYOklrqT+eMYhTrM2+2GBTfU
vPOTZ3Fsp3FZZ0jvP8XL4uiAUF2/VvLxbCP44WkcOG9+PNAVvpac9KKtYnq+kBBT6G0OoKjjRRKc
Uv3iEByI+D8PVJmdnTz1NHZIDHamigC0438bVQBVv4Ar4Wqnp50wIZ6U7FzrKH3l3/EoZGkGXvdZ
kZYpLNHX+zhU2k8iwd4xe3cpFDMxXkIO2kH/3ErBONrK1rayy0EpxSAxgNj2o3hN9eLpfJfByyau
9wixKA1+au0+s/J4nthFZBO6o7EcLujH0XhEeOFUNond6yvHHBOEUfHufY3UTojUDLeG3j9nOF1V
hMPWTa8J3/VG3zjMpQb2t0E0owRRat5O05G8+Rc+DyqNVaKPkRUSfWcxU4w4Lhy8RgkW5ZLBhSXu
d6ozn02Dnf3Gw72un1/6WT67NhbQMcvizZ2b0DS0OMuFJChNOzkAds5XkKWeA0ceUtIJBeAT3Gyd
M9KZdU27PAbRm4hSYmQ0n7HVIL1owBzLkiXq5S/wHI+6i5LJlgFW/E7Nb1rWBm7SM193BFl4J6JH
8SasuBouMb/vFcuT1rcfCfoFovQEkyJBV1eEvOq8Uo6IZEQUFaeTiIfEnyRQ6hbzrHXVUJRZYJ2U
c5lqd79Qv6u7MUSAF3ZnXded5TyccfRvFY9LjcSl3SVMW29XnetQPqw7VBIDdoccKuyUz+xJLarE
b96T4+UBZc4msGsE5sglgBCTavlNKEVnhEX1uqghdMsii0NDEzh9mUN40ZMwgxFKLuxWs4IbKNaf
w85DnjIoC0UerwP8KJPwmFNYohz6z9ourBxWJ6tYP1StGqGOS8QDRj7nBWx+UlhDD0LCUGjd+hvL
mtFow4tUwJ/aqX6grfih4EbGqGGeKcOtEWexliQFTJmGlTIumqpdG1fDaYlrTbFnxUkH18xReFwV
DGYfOvuFPZh4yIz7/YcwQBEtLNKU/B9NV37o7IoQQyIaa1G39Qig9cEAI0zhbF2itmMx92zIWeQO
1DVjrTR5gv3hYszvLZvgYLSY3HqC/JqYFTBsbh2I3N5JXmmIRaViwb2sgs3aG7QtHeoVWz60dvg1
bjqNOiX2X8bbQ4g2/ozrp0lGAwhmiRhRIo2N6IpyCYkxwrZ+3BxUbpZF9ib+cPncpbo0JljKoRSl
VtRtMVrsjUGig0q7OZo2smOWMOp/br1KJKsEAqsRMjtHYzJW3D0TAUfuD0VedXAz65itl+ml15xM
PHSqZbDmzl+flOZaO5BQcikeLZOoM7T0UeFzD6zL0hyln899tf0JaymR93iPwTEiSaA9e73piRtr
XmmRlV3OxV7lapUdDoqd+wi0MbSj652AC6QknJPzqqF5Z6WRyWYIAfwaoWBKeGxJlQZJUYSz0T4o
FkoWHhQsWMoY+ukgkHL3hm49xCxDXqMatl3hvRRmFl0C5SwKrJlyJxHaIeZ8Jqk5DikyKoz474cu
dQ+6z7F6+Bd+uAKejX4CiQz5ZyjaVdUd0uuNjIdlKhjUKsUr2Azp4MbfrEm+7+NT2Au/gQSrhnz5
4Vk6oCNCNRZz00tJcQi7h4oqQeHCvmyI6coSaW0NamYHbcpE0id7fnPnCrrXiXz4+GoX/jZ1Dp1n
WB7YtH01LY2alvgrW8avSSQfy0y9pS0ObhYa37TfiOYOhz6qRsqUJr4epWwR8AyLoTtkafqDcnHB
Y42Pj9DiC+o+GAsz2hVm67Qs6jrlZJv5E5BnR2VmGNs9D3cnb2WA+cd+wQZ4MLxsNKWvdGfLD1S9
/JD13YLjFxF9qVU2gz75K4ityyXfLCtBdM5MrYCWr2G0qNtAR1O2CxLCc4TiuvIqm2Nh3DujA7Ss
yHZ+4AYqGrVBXuCaO356zUZMQC6AexULV86KGTuSpE5liMQoKEfSIwUb6VTqOegMtzX6GiVag+Pz
o8BcE06EjeJWDmU9Vj5YylFYGs/bRsAK0PDJIHPqYeueAZTZru1kFOK0Bvtfv+aQVMlEkwjDEcuX
DiNHKqDYaZra7xWsJAzwioBF7BWeOpiNiWL2JhPYRh2tJceg3k6yLp6SU4Kk7tf/cAmCvhRmbXxB
WFwtNiDMDLT4AkPpFjYphUJInA/mC+16E+uCgT3TvXpFkid1yDf5GI/512vZo/PH3jXkrUbWqbWW
hffg94j+a1d5b49sBS3w2FeWBV6llvniwO6SWe7xAaXDEmek+ir7j35yeX9bzZbdYyb1B5ra9lzd
yb2E4FQ+BFtmfqiCNd4FVg++aVwX3IQE/w63GWHSXsjcThnaI/RzynQuhNCwQtWo9WDCSWplH7nL
DkHjnk/9Qna/230/O96ol78phW246+CL7pywIE7hTEtTdJUZ6ryYHbl7YanUvz14gqecqe/nfB+4
6YQmMDS91ApdhMTvXZSVjlCoKiUt9xbRyDvYyua6bmKrDoBi2oKjPXm6KblhV1YSKLz6FeFdODDK
b+zv7vT9S44XLOyMTS985I5tXtwumhLikDqJMTPkVc29Py2cMNZod7vIsen5pEgt2+oB3ktEC+Os
51zm0oXF4JAgv2MZ6YUXMR6htQ6f3HU7sXRloY0iFaFas74PTa8PxiIgmTo2u2lGdm76asqVVKvj
M3URHDxJlrANsKIvYC1p+9Z4hZRzLq7aEFjAzb/M3h9bTb+4M2A8JDMC59CvCo110WebGc/IIGKz
J9r9+hJ1za2nis4p+3KNZBJsBQt+kFWNUv0W8pLEBe8sWKHntOTcSOn512XrPpmNCNcX/7/dqdUd
IOK3rOTJ3+D48yShybhLtPteUZhSDYblRy+zJSYLGXyo1HHXG4XtAHvfWMLJYn0WXKmM8eH1zb/O
ytFwqVqVvMMCFyWu0sKwNbMTFq3NY52ocU8L4WZ92vSSE5+n9SZoH6Ch/ZPJB5XKpX6jhFJr7D+d
Ig0/1bgKNLPSAph/ff01jDsKKeior7M0AjxdiAMN3ON72wpnD5JkuSTR1RMDtgQqJ33B73qfwUPq
rCkS9yUc/PF/TzDZuRYUHNaEVqna+TW1IbBDBy/L5gDJeYzmjnLZgKg/otPEGeXMoFPypgfV2B4f
+xHCIhjA8cFXlDb3W3CaMkLVUOCP89eTkV2S+t6CVtWdBAADQyw0/NlbviTg7t9ADKvB0ZuXFATR
L0g+V1Ff5Oc0udTrvb8BJBcwM5K9fKwdlZybOnkUfGv1RpNcvfaAxBYPVP2t4p1IfZUXLc1N691X
ocTxDTATu7pXF1WgcBm/fvwEg8PO2p4xOiIwc1c3Wdc4c6OqWW/pjmfh1cnJp/4MBaCHJQU6sJvY
3rQuEgL/7JjGaph/9jd2huGZx/Igo19DkKtLp/JA6O/oa9Hi58wwuivRqX+I2BgUIkdmPNNbmCUC
oWhnIUT35vLJHWSywrPtnyw0Ivm659aw99rmmwsyrAv3gtqm+KTrsQiecY1P9HbguaP/s2B74NNO
5Bf4jBI/aVuV4byNyU8M4JZyIOGBd1meT8u94TnpVlDRzRHGx8NHqr4qoZvybMBaSIjyef6+ed1S
+8+d3Gf9kUdagc4I3JPr435a6K0m3RL5FZ0ngwVgw3/oZsfUlIbXDfjlRS93Lp5X9HUrRIHt/nQl
y2abe8kdeG2+Q7OSfHgy5Q6iiUgNyop2pa/kB6euZmnGUdOJIZToGfRFjarEcroM8g2IVHPydAYG
tOG2ex55Jwz1Go3kPfAN3LjuOqTFMWiPjKvlcgdEUxgSzdkPy3wJnMzbSP7JCg6gCvClLiWkNUNB
Tl+aaPDUn1Z+C9/dgqeHq0KjejmTZP8pYHPzg3QYYbBxUAAjSxgoyi/T7G+Q85G6wQdJIWJJZQ77
iKrOpZNlGZRqYBNmvKHt6YKg2iJSkq0Sdmmi1V4v5ImRnCY0l0VQYGPdbgw0qgk6mo+2rZiVhZ0z
ZWJg32Mp68UcvRRfvupshzxeSwzpIi8cy1JsiE2Z/apRomcTbuRyn4BFSm2b2WS54BJMqhKAhY3I
ggTXK1aqrcuZTMImJT7tyju7Ubu1nKN7aLu18GF7pv+RAPSp1snJ1B3+58wkkFecLG5tms8u8K6R
gG1FEPtV6miWonzLfs2FZwy54luAhwZHOC/WT+i3tbSvmm39+pOxORme5OTHTzEcLQltA1ffgjFR
633OqmIHWAfK5/tuZl6BDa4CahXm1FzHYy5irj58u45q8BanZiHV+kEVevaGbSSJk7rkD8zUI8fO
6i8vfRC8++EqXCn4uZ3TN4ac2fCm7EvxnZg0i56Liv0x0xyxWzPvqJP5bymU++BBIm8Oj7xrOyaZ
uZnZcatLoNkhDSp3tk21lsgyJtAFyZtfH+PLRC5AmEqkmxQk+Bb005Fgau1QWn4G7T4+OKJoCWi8
4ePvh6qB5Gnr3zJSWs9fzKDl3PX/0siTMBqvq0rICURCZSAn25UC/nAbnw79UUzMTm2ZQ1XCqPKU
y8lbpvQ2QdpDjV2ICv3GdrJMGwI1ZiUUm/KodiHUINyQzV1go5Y/owXV8Du4XM7+5IVovj6IZgVi
GmNm1ihGz+Tgnyc/0SD0dYgcdmOG9VEfUz0bSOs6G7L/OkS5cPfs7td4soS/doIsV+o8uutQuZcy
Z+nIjONG7r/dY8EHOHrNdr1n0gHl4HhDgdGAFo8ZRuH+uHFeJKhRTJlDBNtddKnnAwiaWP9s6V/0
hNM0R4XTB+fclhEQQyS7rrXvE6ht8C6M8hEP+pCfGu8RwklUmz9dKhxeSxLRManLmkrdVWj3VvdA
gzkBOprX7hyVEeHX7FR2YxbeSGi+aWqsjhpA3WEBfKIcP/z+GkdaKOUSeCwtK3YPU18wGC8BQM+4
aZveT3b4wAUIEKM7PRV1Md3gIfF8HOsf7nuYkO/s2RxHYiD+7uwjk9RfUWouJhIL8rGvzxoc4alk
XsGJ2y+U0+efd/teSDMbKnOEpl00TWezg038TqNe8mK+DZpIKlWq3SOoEadGKDOXZG/bl6s5LeMk
RtR6aHrbLiHgqwzfNRZihMGLLwdVm2DTuYqO0CUnipFvzyzGYHeE94bJ/V26DRkzrLXlCCdABoCU
HBfvb8sl2gPINIakFo9hvxaPsTbYriYvCqsUZoBUAg7NZifgMpiT91gfHzs0fVXtvP1dwOTjVTxV
wmQujbOSk/wW5rZYQ+PgJTYU6l1oSm1F9zA3DK3c/HZa5+F+HfYErgLsm9yvI4djaqE7ZptgJqYe
JrilufWSf5X407j+K/cIsjlLkhHZFIn7el4yJc2Biwh8gZWl31JIZoh6tSB0UVL3IPyZjHlO/Lir
m+vvcL0OIBUOrfOTMi3vSjOPSHLrNUJm8FDOVPTJmQYY+kBWBaUN72x0GlYOS/lzOxFZQiu8+llf
zFXpFpdQVrCgBlP7DZOigEHxyaOI3klbCgXlvxEZmGmi1R5YbYhZTFqh24yqbxmLJfuYwrVWcivv
ACH9grGQOCrvWTDz9MpNHen5PhXH107oeEg/t3M5R3qDij8zN2aTYe2yqJQ8s9P4P1yuzVN6u9RQ
YaS2BbdNhpshZaN+PQPZprhlLq/xI85xyeSSY/tcw+wcUGzI3zr25BxR3my1TkSUEyUukXzgQc+G
BtWaouj/QeEJi0ges8ZT6nP+W20yzuqmpVj1N2QXK1NQyVLmpNRP8qk25PbCxZuM+B9pNonakqlS
JE9KzFspF5uR36ZxuETEd9LqCpeCdyEQwUSMtAF/nvaii4YPoLIFPbkGfbDXdQYavDIRp1aNC5Wv
WaE2EB7xlp0u8/3oAoM7VLndlePM9y+RjL7WfOOxoN+o1/ZLWHarAC2O8wWb+huSliKN4KQP6riA
Ps3LmHX3B6wAM3wDw2ui9G43ii2IZqKQhrfxeXXfK0d1edF+qCObHYPMZUNgFdOcdY9ulvWdRbSe
8Yu0Chs1jkGXOvnP9p1bFf1m8YyxPnH3zU3MCCbFx907eDsXqq7nSUIFE74Rhuq19K2ejEldgXzf
ZY6Kw92lQlXnRBSPBt13HPoPhQrielsQ0b/PYzbYNB/Hn7ScrnGQ63wi/cvbKdQ7jJXDAAQZTD5w
FY001pdgJSQQNbQNHhuMXeP8DYtE+GFeXZ3CLlvERIGu+mW8mPMYGmtYPZPSjdleTG9duJ/z4O74
gHUp7iCyQOIojPhNYPZKt+P8+sh3ufjuvzSUdjhIImrwNUhz5X951iKb2weg2jai6JeYh2XrK76j
vRTGOHJ5CGfNvII6W1x8dIj3jeZcq3Werf3Ch44iyaKPias+7p5hg720QItDL7tQD0/Aa8B50TfV
2hqNGxBVwa6c6SM0uOdelIJYiJcW3Z7+zS5fblraBPlEpv+FQT3XfjIHcxHBQml3TmS3bbAsxSi0
jdI6kRdYTNJ7+395Dt85hScWKAOwuV28BCKvHKAAayWO8dPkHlm5tV09iF+SDI9QSlP27NIQvB/O
eXZgkuGzEHRVUxBnS5O/vk/P7b/4BoJMPOMRkZ3N61W/vBdzudL9kXuhK82Ij0UtGAkgOgbBIZg6
GsRuBajtgJgmMKzNr8PCQVX8BYn3lMMGOeySoTS+AudhUeku1F9uWSx4EQMC3ZqYlv+Ut5JLKGi/
jHXtbp+MiHhNyft0/axE9nbXXruAEFsC5yXtQeTZWq1An89/VGznYG6y+Gju8zZ23neSpIxtNmi/
JyCE6/8OpkTKZ0zht4IbHxPW2rQJNb3Ys4T6VMwoTsa0e8vm77SAyLOolDKf/ed1fRmxCVz2dEW+
4A11jnwNuVVXr4uuFmLVF6vwzRu+v8LoslgnRGfFbEDEApzRISb7MPid3oBD89jhbVC6OdvDplp7
sG0YCdnfy8lsYw1RhOfq7gtyNmOxVWl+itrj05+gw7UURk14bzXAdEyY+Q3zph1jZz6tmFKJ4S2x
moofyj5HBqK/uYRmo67oQEJz6C5xSgBhGtzdHxFZQZCxOybpGI/jfyAHPqPKr2QvfVpIXho+oDa1
h5ZpKG0bd92ezy8T8FyML9cYWG4dMkxoMCQ9I62tnz1aLX5gi/tHzANraU0uTTqMGt8RqeR7lZUC
crZV/zsdxvdxEc/1nygNOt0X4Hork+2XyJUzT2xycyFeKuFqLaNH5TWsXHDtKKZQA9rHyQswRpYi
g9ChQQ9Uts7BOsPoHphQ1svPZQmcSYhetlkHj7N1yaHMLPcxois+fJ1yjOqNj9q0QNpHlDPpW+Hu
1nc/UXqBkegOExeKUfo2FqyFIng7g15YwiM3mUZptizqwA48O8+k7ionKh4xPow3vpDwIS8uxfPM
Vx2/drmzK2FSkWskZavZLVuEX1ry2StWVrozQgb1HEAerst5bWbZviM794wCyLax1+wDq7s985xJ
+ayzOi1c/EnbcVu7sQ3TXPj5+JfwE0Te6bB0B+mU/BYkQG8QMr7kMDwFV1KAlBTu+SeIk4abbJVx
46FMydlg/ii/ruKlSAATUuxuHWWoq7EG1n9PbiuXSDR/msxfaZNFJgYRjCdMZHOt6u3JPzJPpdmA
Nbev0ggFARMR6JOxPSN147+iyiYrV5FTF1CUKnkbGHF4tQijgqn6OFj4TXWtsqwuNbmCvGuu5PVH
akprZf5QBtmaJIO1jaY21PNTWTqs+2NiGEdC1srxo6W8CpS/J2NvR4gV/tDI5dlziFWdwSjG6Dmz
tfd1SSlwrgN9UzdVDE6JBUEVk0ZtBazTDosYzXe3WvySbj6WFUW9vRJ1UDPVl8+in8JGxLGcxqtr
D1NaNW808jy0YTl0HQX5/8Na+BLvax/ZT2CVnomVEhA6HvCX6aD0Ysw5r29NZR8DdRFm2/UTcm3o
bFtILQDy7+/zKKGtdErRkAcfFciQxYfnPi0GY+7pL2gQnaz0L5n0/sd8BswXLsIXqv8ex2hJ4sR7
TLZekMYo8EHa4yU76ehgADQkXeBnkRqqQw==
`protect end_protected
